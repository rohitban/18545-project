

module pwm_thresh_96k
    (input  logic [9:0] mult_val,
     output logic [10:0] pwm_thresh);

    always_comb begin
        case(mult_val)
            10'h0: pwm_thresh = 11'd0;
            10'h1: pwm_thresh = 11'd1;
            10'h2: pwm_thresh = 11'd2;
            10'h3: pwm_thresh = 11'd3;
            10'h4: pwm_thresh = 11'd4;
            10'h5: pwm_thresh = 11'd5;
            10'h6: pwm_thresh = 11'd6;
            10'h7: pwm_thresh = 11'd7;
            10'h8: pwm_thresh = 11'd8;
            10'h9: pwm_thresh = 11'd9;
            10'ha: pwm_thresh = 11'd10;
            10'hb: pwm_thresh = 11'd11;
            10'hc: pwm_thresh = 11'd12;
            10'hd: pwm_thresh = 11'd13;
            10'he: pwm_thresh = 11'd14;
            10'hf: pwm_thresh = 11'd15;
            10'h10: pwm_thresh = 11'd16;
            10'h11: pwm_thresh = 11'd17;
            10'h12: pwm_thresh = 11'd18;
            10'h13: pwm_thresh = 11'd19;
            10'h14: pwm_thresh = 11'd20;
            10'h15: pwm_thresh = 11'd21;
            10'h16: pwm_thresh = 11'd22;
            10'h17: pwm_thresh = 11'd23;
            10'h18: pwm_thresh = 11'd24;
            10'h19: pwm_thresh = 11'd25;
            10'h1a: pwm_thresh = 11'd26;
            10'h1b: pwm_thresh = 11'd27;
            10'h1c: pwm_thresh = 11'd28;
            10'h1d: pwm_thresh = 11'd29;
            10'h1e: pwm_thresh = 11'd30;
            10'h1f: pwm_thresh = 11'd31;
            10'h20: pwm_thresh = 11'd32;
            10'h21: pwm_thresh = 11'd33;
            10'h22: pwm_thresh = 11'd34;
            10'h23: pwm_thresh = 11'd35;
            10'h24: pwm_thresh = 11'd36;
            10'h25: pwm_thresh = 11'd37;
            10'h26: pwm_thresh = 11'd38;
            10'h27: pwm_thresh = 11'd39;
            10'h28: pwm_thresh = 11'd40;
            10'h29: pwm_thresh = 11'd41;
            10'h2a: pwm_thresh = 11'd42;
            10'h2b: pwm_thresh = 11'd43;
            10'h2c: pwm_thresh = 11'd44;
            10'h2d: pwm_thresh = 11'd45;
            10'h2e: pwm_thresh = 11'd46;
            10'h2f: pwm_thresh = 11'd47;
            10'h30: pwm_thresh = 11'd48;
            10'h31: pwm_thresh = 11'd49;
            10'h32: pwm_thresh = 11'd50;
            10'h33: pwm_thresh = 11'd51;
            10'h34: pwm_thresh = 11'd52;
            10'h35: pwm_thresh = 11'd53;
            10'h36: pwm_thresh = 11'd55;
            10'h37: pwm_thresh = 11'd56;
            10'h38: pwm_thresh = 11'd57;
            10'h39: pwm_thresh = 11'd58;
            10'h3a: pwm_thresh = 11'd59;
            10'h3b: pwm_thresh = 11'd60;
            10'h3c: pwm_thresh = 11'd61;
            10'h3d: pwm_thresh = 11'd62;
            10'h3e: pwm_thresh = 11'd63;
            10'h3f: pwm_thresh = 11'd64;
            10'h40: pwm_thresh = 11'd65;
            10'h41: pwm_thresh = 11'd66;
            10'h42: pwm_thresh = 11'd67;
            10'h43: pwm_thresh = 11'd68;
            10'h44: pwm_thresh = 11'd69;
            10'h45: pwm_thresh = 11'd70;
            10'h46: pwm_thresh = 11'd71;
            10'h47: pwm_thresh = 11'd72;
            10'h48: pwm_thresh = 11'd73;
            10'h49: pwm_thresh = 11'd74;
            10'h4a: pwm_thresh = 11'd75;
            10'h4b: pwm_thresh = 11'd76;
            10'h4c: pwm_thresh = 11'd77;
            10'h4d: pwm_thresh = 11'd78;
            10'h4e: pwm_thresh = 11'd79;
            10'h4f: pwm_thresh = 11'd80;
            10'h50: pwm_thresh = 11'd81;
            10'h51: pwm_thresh = 11'd82;
            10'h52: pwm_thresh = 11'd83;
            10'h53: pwm_thresh = 11'd84;
            10'h54: pwm_thresh = 11'd85;
            10'h55: pwm_thresh = 11'd86;
            10'h56: pwm_thresh = 11'd87;
            10'h57: pwm_thresh = 11'd88;
            10'h58: pwm_thresh = 11'd89;
            10'h59: pwm_thresh = 11'd90;
            10'h5a: pwm_thresh = 11'd91;
            10'h5b: pwm_thresh = 11'd92;
            10'h5c: pwm_thresh = 11'd93;
            10'h5d: pwm_thresh = 11'd94;
            10'h5e: pwm_thresh = 11'd95;
            10'h5f: pwm_thresh = 11'd96;
            10'h60: pwm_thresh = 11'd97;
            10'h61: pwm_thresh = 11'd98;
            10'h62: pwm_thresh = 11'd99;
            10'h63: pwm_thresh = 11'd100;
            10'h64: pwm_thresh = 11'd101;
            10'h65: pwm_thresh = 11'd102;
            10'h66: pwm_thresh = 11'd103;
            10'h67: pwm_thresh = 11'd104;
            10'h68: pwm_thresh = 11'd105;
            10'h69: pwm_thresh = 11'd106;
            10'h6a: pwm_thresh = 11'd107;
            10'h6b: pwm_thresh = 11'd108;
            10'h6c: pwm_thresh = 11'd110;
            10'h6d: pwm_thresh = 11'd111;
            10'h6e: pwm_thresh = 11'd112;
            10'h6f: pwm_thresh = 11'd113;
            10'h70: pwm_thresh = 11'd114;
            10'h71: pwm_thresh = 11'd115;
            10'h72: pwm_thresh = 11'd116;
            10'h73: pwm_thresh = 11'd117;
            10'h74: pwm_thresh = 11'd118;
            10'h75: pwm_thresh = 11'd119;
            10'h76: pwm_thresh = 11'd120;
            10'h77: pwm_thresh = 11'd121;
            10'h78: pwm_thresh = 11'd122;
            10'h79: pwm_thresh = 11'd123;
            10'h7a: pwm_thresh = 11'd124;
            10'h7b: pwm_thresh = 11'd125;
            10'h7c: pwm_thresh = 11'd126;
            10'h7d: pwm_thresh = 11'd127;
            10'h7e: pwm_thresh = 11'd128;
            10'h7f: pwm_thresh = 11'd129;
            10'h80: pwm_thresh = 11'd130;
            10'h81: pwm_thresh = 11'd131;
            10'h82: pwm_thresh = 11'd132;
            10'h83: pwm_thresh = 11'd133;
            10'h84: pwm_thresh = 11'd134;
            10'h85: pwm_thresh = 11'd135;
            10'h86: pwm_thresh = 11'd136;
            10'h87: pwm_thresh = 11'd137;
            10'h88: pwm_thresh = 11'd138;
            10'h89: pwm_thresh = 11'd139;
            10'h8a: pwm_thresh = 11'd140;
            10'h8b: pwm_thresh = 11'd141;
            10'h8c: pwm_thresh = 11'd142;
            10'h8d: pwm_thresh = 11'd143;
            10'h8e: pwm_thresh = 11'd144;
            10'h8f: pwm_thresh = 11'd145;
            10'h90: pwm_thresh = 11'd146;
            10'h91: pwm_thresh = 11'd147;
            10'h92: pwm_thresh = 11'd148;
            10'h93: pwm_thresh = 11'd149;
            10'h94: pwm_thresh = 11'd150;
            10'h95: pwm_thresh = 11'd151;
            10'h96: pwm_thresh = 11'd152;
            10'h97: pwm_thresh = 11'd153;
            10'h98: pwm_thresh = 11'd154;
            10'h99: pwm_thresh = 11'd155;
            10'h9a: pwm_thresh = 11'd156;
            10'h9b: pwm_thresh = 11'd157;
            10'h9c: pwm_thresh = 11'd158;
            10'h9d: pwm_thresh = 11'd159;
            10'h9e: pwm_thresh = 11'd160;
            10'h9f: pwm_thresh = 11'd161;
            10'ha0: pwm_thresh = 11'd162;
            10'ha1: pwm_thresh = 11'd163;
            10'ha2: pwm_thresh = 11'd165;
            10'ha3: pwm_thresh = 11'd166;
            10'ha4: pwm_thresh = 11'd167;
            10'ha5: pwm_thresh = 11'd168;
            10'ha6: pwm_thresh = 11'd169;
            10'ha7: pwm_thresh = 11'd170;
            10'ha8: pwm_thresh = 11'd171;
            10'ha9: pwm_thresh = 11'd172;
            10'haa: pwm_thresh = 11'd173;
            10'hab: pwm_thresh = 11'd174;
            10'hac: pwm_thresh = 11'd175;
            10'had: pwm_thresh = 11'd176;
            10'hae: pwm_thresh = 11'd177;
            10'haf: pwm_thresh = 11'd178;
            10'hb0: pwm_thresh = 11'd179;
            10'hb1: pwm_thresh = 11'd180;
            10'hb2: pwm_thresh = 11'd181;
            10'hb3: pwm_thresh = 11'd182;
            10'hb4: pwm_thresh = 11'd183;
            10'hb5: pwm_thresh = 11'd184;
            10'hb6: pwm_thresh = 11'd185;
            10'hb7: pwm_thresh = 11'd186;
            10'hb8: pwm_thresh = 11'd187;
            10'hb9: pwm_thresh = 11'd188;
            10'hba: pwm_thresh = 11'd189;
            10'hbb: pwm_thresh = 11'd190;
            10'hbc: pwm_thresh = 11'd191;
            10'hbd: pwm_thresh = 11'd192;
            10'hbe: pwm_thresh = 11'd193;
            10'hbf: pwm_thresh = 11'd194;
            10'hc0: pwm_thresh = 11'd195;
            10'hc1: pwm_thresh = 11'd196;
            10'hc2: pwm_thresh = 11'd197;
            10'hc3: pwm_thresh = 11'd198;
            10'hc4: pwm_thresh = 11'd199;
            10'hc5: pwm_thresh = 11'd200;
            10'hc6: pwm_thresh = 11'd201;
            10'hc7: pwm_thresh = 11'd202;
            10'hc8: pwm_thresh = 11'd203;
            10'hc9: pwm_thresh = 11'd204;
            10'hca: pwm_thresh = 11'd205;
            10'hcb: pwm_thresh = 11'd206;
            10'hcc: pwm_thresh = 11'd207;
            10'hcd: pwm_thresh = 11'd208;
            10'hce: pwm_thresh = 11'd209;
            10'hcf: pwm_thresh = 11'd210;
            10'hd0: pwm_thresh = 11'd211;
            10'hd1: pwm_thresh = 11'd212;
            10'hd2: pwm_thresh = 11'd213;
            10'hd3: pwm_thresh = 11'd214;
            10'hd4: pwm_thresh = 11'd215;
            10'hd5: pwm_thresh = 11'd216;
            10'hd6: pwm_thresh = 11'd217;
            10'hd7: pwm_thresh = 11'd218;
            10'hd8: pwm_thresh = 11'd220;
            10'hd9: pwm_thresh = 11'd221;
            10'hda: pwm_thresh = 11'd222;
            10'hdb: pwm_thresh = 11'd223;
            10'hdc: pwm_thresh = 11'd224;
            10'hdd: pwm_thresh = 11'd225;
            10'hde: pwm_thresh = 11'd226;
            10'hdf: pwm_thresh = 11'd227;
            10'he0: pwm_thresh = 11'd228;
            10'he1: pwm_thresh = 11'd229;
            10'he2: pwm_thresh = 11'd230;
            10'he3: pwm_thresh = 11'd231;
            10'he4: pwm_thresh = 11'd232;
            10'he5: pwm_thresh = 11'd233;
            10'he6: pwm_thresh = 11'd234;
            10'he7: pwm_thresh = 11'd235;
            10'he8: pwm_thresh = 11'd236;
            10'he9: pwm_thresh = 11'd237;
            10'hea: pwm_thresh = 11'd238;
            10'heb: pwm_thresh = 11'd239;
            10'hec: pwm_thresh = 11'd240;
            10'hed: pwm_thresh = 11'd241;
            10'hee: pwm_thresh = 11'd242;
            10'hef: pwm_thresh = 11'd243;
            10'hf0: pwm_thresh = 11'd244;
            10'hf1: pwm_thresh = 11'd245;
            10'hf2: pwm_thresh = 11'd246;
            10'hf3: pwm_thresh = 11'd247;
            10'hf4: pwm_thresh = 11'd248;
            10'hf5: pwm_thresh = 11'd249;
            10'hf6: pwm_thresh = 11'd250;
            10'hf7: pwm_thresh = 11'd251;
            10'hf8: pwm_thresh = 11'd252;
            10'hf9: pwm_thresh = 11'd253;
            10'hfa: pwm_thresh = 11'd254;
            10'hfb: pwm_thresh = 11'd255;
            10'hfc: pwm_thresh = 11'd256;
            10'hfd: pwm_thresh = 11'd257;
            10'hfe: pwm_thresh = 11'd258;
            10'hff: pwm_thresh = 11'd259;
            10'h100: pwm_thresh = 11'd260;
            10'h101: pwm_thresh = 11'd261;
            10'h102: pwm_thresh = 11'd262;
            10'h103: pwm_thresh = 11'd263;
            10'h104: pwm_thresh = 11'd264;
            10'h105: pwm_thresh = 11'd265;
            10'h106: pwm_thresh = 11'd266;
            10'h107: pwm_thresh = 11'd267;
            10'h108: pwm_thresh = 11'd268;
            10'h109: pwm_thresh = 11'd269;
            10'h10a: pwm_thresh = 11'd270;
            10'h10b: pwm_thresh = 11'd271;
            10'h10c: pwm_thresh = 11'd272;
            10'h10d: pwm_thresh = 11'd273;
            10'h10e: pwm_thresh = 11'd275;
            10'h10f: pwm_thresh = 11'd276;
            10'h110: pwm_thresh = 11'd277;
            10'h111: pwm_thresh = 11'd278;
            10'h112: pwm_thresh = 11'd279;
            10'h113: pwm_thresh = 11'd280;
            10'h114: pwm_thresh = 11'd281;
            10'h115: pwm_thresh = 11'd282;
            10'h116: pwm_thresh = 11'd283;
            10'h117: pwm_thresh = 11'd284;
            10'h118: pwm_thresh = 11'd285;
            10'h119: pwm_thresh = 11'd286;
            10'h11a: pwm_thresh = 11'd287;
            10'h11b: pwm_thresh = 11'd288;
            10'h11c: pwm_thresh = 11'd289;
            10'h11d: pwm_thresh = 11'd290;
            10'h11e: pwm_thresh = 11'd291;
            10'h11f: pwm_thresh = 11'd292;
            10'h120: pwm_thresh = 11'd293;
            10'h121: pwm_thresh = 11'd294;
            10'h122: pwm_thresh = 11'd295;
            10'h123: pwm_thresh = 11'd296;
            10'h124: pwm_thresh = 11'd297;
            10'h125: pwm_thresh = 11'd298;
            10'h126: pwm_thresh = 11'd299;
            10'h127: pwm_thresh = 11'd300;
            10'h128: pwm_thresh = 11'd301;
            10'h129: pwm_thresh = 11'd302;
            10'h12a: pwm_thresh = 11'd303;
            10'h12b: pwm_thresh = 11'd304;
            10'h12c: pwm_thresh = 11'd305;
            10'h12d: pwm_thresh = 11'd306;
            10'h12e: pwm_thresh = 11'd307;
            10'h12f: pwm_thresh = 11'd308;
            10'h130: pwm_thresh = 11'd309;
            10'h131: pwm_thresh = 11'd310;
            10'h132: pwm_thresh = 11'd311;
            10'h133: pwm_thresh = 11'd312;
            10'h134: pwm_thresh = 11'd313;
            10'h135: pwm_thresh = 11'd314;
            10'h136: pwm_thresh = 11'd315;
            10'h137: pwm_thresh = 11'd316;
            10'h138: pwm_thresh = 11'd317;
            10'h139: pwm_thresh = 11'd318;
            10'h13a: pwm_thresh = 11'd319;
            10'h13b: pwm_thresh = 11'd320;
            10'h13c: pwm_thresh = 11'd321;
            10'h13d: pwm_thresh = 11'd322;
            10'h13e: pwm_thresh = 11'd323;
            10'h13f: pwm_thresh = 11'd324;
            10'h140: pwm_thresh = 11'd325;
            10'h141: pwm_thresh = 11'd326;
            10'h142: pwm_thresh = 11'd327;
            10'h143: pwm_thresh = 11'd328;
            10'h144: pwm_thresh = 11'd330;
            10'h145: pwm_thresh = 11'd331;
            10'h146: pwm_thresh = 11'd332;
            10'h147: pwm_thresh = 11'd333;
            10'h148: pwm_thresh = 11'd334;
            10'h149: pwm_thresh = 11'd335;
            10'h14a: pwm_thresh = 11'd336;
            10'h14b: pwm_thresh = 11'd337;
            10'h14c: pwm_thresh = 11'd338;
            10'h14d: pwm_thresh = 11'd339;
            10'h14e: pwm_thresh = 11'd340;
            10'h14f: pwm_thresh = 11'd341;
            10'h150: pwm_thresh = 11'd342;
            10'h151: pwm_thresh = 11'd343;
            10'h152: pwm_thresh = 11'd344;
            10'h153: pwm_thresh = 11'd345;
            10'h154: pwm_thresh = 11'd346;
            10'h155: pwm_thresh = 11'd347;
            10'h156: pwm_thresh = 11'd348;
            10'h157: pwm_thresh = 11'd349;
            10'h158: pwm_thresh = 11'd350;
            10'h159: pwm_thresh = 11'd351;
            10'h15a: pwm_thresh = 11'd352;
            10'h15b: pwm_thresh = 11'd353;
            10'h15c: pwm_thresh = 11'd354;
            10'h15d: pwm_thresh = 11'd355;
            10'h15e: pwm_thresh = 11'd356;
            10'h15f: pwm_thresh = 11'd357;
            10'h160: pwm_thresh = 11'd358;
            10'h161: pwm_thresh = 11'd359;
            10'h162: pwm_thresh = 11'd360;
            10'h163: pwm_thresh = 11'd361;
            10'h164: pwm_thresh = 11'd362;
            10'h165: pwm_thresh = 11'd363;
            10'h166: pwm_thresh = 11'd364;
            10'h167: pwm_thresh = 11'd365;
            10'h168: pwm_thresh = 11'd366;
            10'h169: pwm_thresh = 11'd367;
            10'h16a: pwm_thresh = 11'd368;
            10'h16b: pwm_thresh = 11'd369;
            10'h16c: pwm_thresh = 11'd370;
            10'h16d: pwm_thresh = 11'd371;
            10'h16e: pwm_thresh = 11'd372;
            10'h16f: pwm_thresh = 11'd373;
            10'h170: pwm_thresh = 11'd374;
            10'h171: pwm_thresh = 11'd375;
            10'h172: pwm_thresh = 11'd376;
            10'h173: pwm_thresh = 11'd377;
            10'h174: pwm_thresh = 11'd378;
            10'h175: pwm_thresh = 11'd379;
            10'h176: pwm_thresh = 11'd380;
            10'h177: pwm_thresh = 11'd381;
            10'h178: pwm_thresh = 11'd382;
            10'h179: pwm_thresh = 11'd384;
            10'h17a: pwm_thresh = 11'd385;
            10'h17b: pwm_thresh = 11'd386;
            10'h17c: pwm_thresh = 11'd387;
            10'h17d: pwm_thresh = 11'd388;
            10'h17e: pwm_thresh = 11'd389;
            10'h17f: pwm_thresh = 11'd390;
            10'h180: pwm_thresh = 11'd391;
            10'h181: pwm_thresh = 11'd392;
            10'h182: pwm_thresh = 11'd393;
            10'h183: pwm_thresh = 11'd394;
            10'h184: pwm_thresh = 11'd395;
            10'h185: pwm_thresh = 11'd396;
            10'h186: pwm_thresh = 11'd397;
            10'h187: pwm_thresh = 11'd398;
            10'h188: pwm_thresh = 11'd399;
            10'h189: pwm_thresh = 11'd400;
            10'h18a: pwm_thresh = 11'd401;
            10'h18b: pwm_thresh = 11'd402;
            10'h18c: pwm_thresh = 11'd403;
            10'h18d: pwm_thresh = 11'd404;
            10'h18e: pwm_thresh = 11'd405;
            10'h18f: pwm_thresh = 11'd406;
            10'h190: pwm_thresh = 11'd407;
            10'h191: pwm_thresh = 11'd408;
            10'h192: pwm_thresh = 11'd409;
            10'h193: pwm_thresh = 11'd410;
            10'h194: pwm_thresh = 11'd411;
            10'h195: pwm_thresh = 11'd412;
            10'h196: pwm_thresh = 11'd413;
            10'h197: pwm_thresh = 11'd414;
            10'h198: pwm_thresh = 11'd415;
            10'h199: pwm_thresh = 11'd416;
            10'h19a: pwm_thresh = 11'd417;
            10'h19b: pwm_thresh = 11'd418;
            10'h19c: pwm_thresh = 11'd419;
            10'h19d: pwm_thresh = 11'd420;
            10'h19e: pwm_thresh = 11'd421;
            10'h19f: pwm_thresh = 11'd422;
            10'h1a0: pwm_thresh = 11'd423;
            10'h1a1: pwm_thresh = 11'd424;
            10'h1a2: pwm_thresh = 11'd425;
            10'h1a3: pwm_thresh = 11'd426;
            10'h1a4: pwm_thresh = 11'd427;
            10'h1a5: pwm_thresh = 11'd428;
            10'h1a6: pwm_thresh = 11'd429;
            10'h1a7: pwm_thresh = 11'd430;
            10'h1a8: pwm_thresh = 11'd431;
            10'h1a9: pwm_thresh = 11'd432;
            10'h1aa: pwm_thresh = 11'd433;
            10'h1ab: pwm_thresh = 11'd434;
            10'h1ac: pwm_thresh = 11'd435;
            10'h1ad: pwm_thresh = 11'd436;
            10'h1ae: pwm_thresh = 11'd437;
            10'h1af: pwm_thresh = 11'd439;
            10'h1b0: pwm_thresh = 11'd440;
            10'h1b1: pwm_thresh = 11'd441;
            10'h1b2: pwm_thresh = 11'd442;
            10'h1b3: pwm_thresh = 11'd443;
            10'h1b4: pwm_thresh = 11'd444;
            10'h1b5: pwm_thresh = 11'd445;
            10'h1b6: pwm_thresh = 11'd446;
            10'h1b7: pwm_thresh = 11'd447;
            10'h1b8: pwm_thresh = 11'd448;
            10'h1b9: pwm_thresh = 11'd449;
            10'h1ba: pwm_thresh = 11'd450;
            10'h1bb: pwm_thresh = 11'd451;
            10'h1bc: pwm_thresh = 11'd452;
            10'h1bd: pwm_thresh = 11'd453;
            10'h1be: pwm_thresh = 11'd454;
            10'h1bf: pwm_thresh = 11'd455;
            10'h1c0: pwm_thresh = 11'd456;
            10'h1c1: pwm_thresh = 11'd457;
            10'h1c2: pwm_thresh = 11'd458;
            10'h1c3: pwm_thresh = 11'd459;
            10'h1c4: pwm_thresh = 11'd460;
            10'h1c5: pwm_thresh = 11'd461;
            10'h1c6: pwm_thresh = 11'd462;
            10'h1c7: pwm_thresh = 11'd463;
            10'h1c8: pwm_thresh = 11'd464;
            10'h1c9: pwm_thresh = 11'd465;
            10'h1ca: pwm_thresh = 11'd466;
            10'h1cb: pwm_thresh = 11'd467;
            10'h1cc: pwm_thresh = 11'd468;
            10'h1cd: pwm_thresh = 11'd469;
            10'h1ce: pwm_thresh = 11'd470;
            10'h1cf: pwm_thresh = 11'd471;
            10'h1d0: pwm_thresh = 11'd472;
            10'h1d1: pwm_thresh = 11'd473;
            10'h1d2: pwm_thresh = 11'd474;
            10'h1d3: pwm_thresh = 11'd475;
            10'h1d4: pwm_thresh = 11'd476;
            10'h1d5: pwm_thresh = 11'd477;
            10'h1d6: pwm_thresh = 11'd478;
            10'h1d7: pwm_thresh = 11'd479;
            10'h1d8: pwm_thresh = 11'd480;
            10'h1d9: pwm_thresh = 11'd481;
            10'h1da: pwm_thresh = 11'd482;
            10'h1db: pwm_thresh = 11'd483;
            10'h1dc: pwm_thresh = 11'd484;
            10'h1dd: pwm_thresh = 11'd485;
            10'h1de: pwm_thresh = 11'd486;
            10'h1df: pwm_thresh = 11'd487;
            10'h1e0: pwm_thresh = 11'd488;
            10'h1e1: pwm_thresh = 11'd489;
            10'h1e2: pwm_thresh = 11'd490;
            10'h1e3: pwm_thresh = 11'd491;
            10'h1e4: pwm_thresh = 11'd492;
            10'h1e5: pwm_thresh = 11'd494;
            10'h1e6: pwm_thresh = 11'd495;
            10'h1e7: pwm_thresh = 11'd496;
            10'h1e8: pwm_thresh = 11'd497;
            10'h1e9: pwm_thresh = 11'd498;
            10'h1ea: pwm_thresh = 11'd499;
            10'h1eb: pwm_thresh = 11'd500;
            10'h1ec: pwm_thresh = 11'd501;
            10'h1ed: pwm_thresh = 11'd502;
            10'h1ee: pwm_thresh = 11'd503;
            10'h1ef: pwm_thresh = 11'd504;
            10'h1f0: pwm_thresh = 11'd505;
            10'h1f1: pwm_thresh = 11'd506;
            10'h1f2: pwm_thresh = 11'd507;
            10'h1f3: pwm_thresh = 11'd508;
            10'h1f4: pwm_thresh = 11'd509;
            10'h1f5: pwm_thresh = 11'd510;
            10'h1f6: pwm_thresh = 11'd511;
            10'h1f7: pwm_thresh = 11'd512;
            10'h1f8: pwm_thresh = 11'd513;
            10'h1f9: pwm_thresh = 11'd514;
            10'h1fa: pwm_thresh = 11'd515;
            10'h1fb: pwm_thresh = 11'd516;
            10'h1fc: pwm_thresh = 11'd517;
            10'h1fd: pwm_thresh = 11'd518;
            10'h1fe: pwm_thresh = 11'd519;
            10'h1ff: pwm_thresh = 11'd520;
            10'h200: pwm_thresh = 11'd521;
            10'h201: pwm_thresh = 11'd522;
            10'h202: pwm_thresh = 11'd523;
            10'h203: pwm_thresh = 11'd524;
            10'h204: pwm_thresh = 11'd525;
            10'h205: pwm_thresh = 11'd526;
            10'h206: pwm_thresh = 11'd527;
            10'h207: pwm_thresh = 11'd528;
            10'h208: pwm_thresh = 11'd529;
            10'h209: pwm_thresh = 11'd530;
            10'h20a: pwm_thresh = 11'd531;
            10'h20b: pwm_thresh = 11'd532;
            10'h20c: pwm_thresh = 11'd533;
            10'h20d: pwm_thresh = 11'd534;
            10'h20e: pwm_thresh = 11'd535;
            10'h20f: pwm_thresh = 11'd536;
            10'h210: pwm_thresh = 11'd537;
            10'h211: pwm_thresh = 11'd538;
            10'h212: pwm_thresh = 11'd539;
            10'h213: pwm_thresh = 11'd540;
            10'h214: pwm_thresh = 11'd541;
            10'h215: pwm_thresh = 11'd542;
            10'h216: pwm_thresh = 11'd543;
            10'h217: pwm_thresh = 11'd544;
            10'h218: pwm_thresh = 11'd545;
            10'h219: pwm_thresh = 11'd546;
            10'h21a: pwm_thresh = 11'd547;
            10'h21b: pwm_thresh = 11'd549;
            10'h21c: pwm_thresh = 11'd550;
            10'h21d: pwm_thresh = 11'd551;
            10'h21e: pwm_thresh = 11'd552;
            10'h21f: pwm_thresh = 11'd553;
            10'h220: pwm_thresh = 11'd554;
            10'h221: pwm_thresh = 11'd555;
            10'h222: pwm_thresh = 11'd556;
            10'h223: pwm_thresh = 11'd557;
            10'h224: pwm_thresh = 11'd558;
            10'h225: pwm_thresh = 11'd559;
            10'h226: pwm_thresh = 11'd560;
            10'h227: pwm_thresh = 11'd561;
            10'h228: pwm_thresh = 11'd562;
            10'h229: pwm_thresh = 11'd563;
            10'h22a: pwm_thresh = 11'd564;
            10'h22b: pwm_thresh = 11'd565;
            10'h22c: pwm_thresh = 11'd566;
            10'h22d: pwm_thresh = 11'd567;
            10'h22e: pwm_thresh = 11'd568;
            10'h22f: pwm_thresh = 11'd569;
            10'h230: pwm_thresh = 11'd570;
            10'h231: pwm_thresh = 11'd571;
            10'h232: pwm_thresh = 11'd572;
            10'h233: pwm_thresh = 11'd573;
            10'h234: pwm_thresh = 11'd574;
            10'h235: pwm_thresh = 11'd575;
            10'h236: pwm_thresh = 11'd576;
            10'h237: pwm_thresh = 11'd577;
            10'h238: pwm_thresh = 11'd578;
            10'h239: pwm_thresh = 11'd579;
            10'h23a: pwm_thresh = 11'd580;
            10'h23b: pwm_thresh = 11'd581;
            10'h23c: pwm_thresh = 11'd582;
            10'h23d: pwm_thresh = 11'd583;
            10'h23e: pwm_thresh = 11'd584;
            10'h23f: pwm_thresh = 11'd585;
            10'h240: pwm_thresh = 11'd586;
            10'h241: pwm_thresh = 11'd587;
            10'h242: pwm_thresh = 11'd588;
            10'h243: pwm_thresh = 11'd589;
            10'h244: pwm_thresh = 11'd590;
            10'h245: pwm_thresh = 11'd591;
            10'h246: pwm_thresh = 11'd592;
            10'h247: pwm_thresh = 11'd593;
            10'h248: pwm_thresh = 11'd594;
            10'h249: pwm_thresh = 11'd595;
            10'h24a: pwm_thresh = 11'd596;
            10'h24b: pwm_thresh = 11'd597;
            10'h24c: pwm_thresh = 11'd598;
            10'h24d: pwm_thresh = 11'd599;
            10'h24e: pwm_thresh = 11'd600;
            10'h24f: pwm_thresh = 11'd601;
            10'h250: pwm_thresh = 11'd602;
            10'h251: pwm_thresh = 11'd604;
            10'h252: pwm_thresh = 11'd605;
            10'h253: pwm_thresh = 11'd606;
            10'h254: pwm_thresh = 11'd607;
            10'h255: pwm_thresh = 11'd608;
            10'h256: pwm_thresh = 11'd609;
            10'h257: pwm_thresh = 11'd610;
            10'h258: pwm_thresh = 11'd611;
            10'h259: pwm_thresh = 11'd612;
            10'h25a: pwm_thresh = 11'd613;
            10'h25b: pwm_thresh = 11'd614;
            10'h25c: pwm_thresh = 11'd615;
            10'h25d: pwm_thresh = 11'd616;
            10'h25e: pwm_thresh = 11'd617;
            10'h25f: pwm_thresh = 11'd618;
            10'h260: pwm_thresh = 11'd619;
            10'h261: pwm_thresh = 11'd620;
            10'h262: pwm_thresh = 11'd621;
            10'h263: pwm_thresh = 11'd622;
            10'h264: pwm_thresh = 11'd623;
            10'h265: pwm_thresh = 11'd624;
            10'h266: pwm_thresh = 11'd625;
            10'h267: pwm_thresh = 11'd626;
            10'h268: pwm_thresh = 11'd627;
            10'h269: pwm_thresh = 11'd628;
            10'h26a: pwm_thresh = 11'd629;
            10'h26b: pwm_thresh = 11'd630;
            10'h26c: pwm_thresh = 11'd631;
            10'h26d: pwm_thresh = 11'd632;
            10'h26e: pwm_thresh = 11'd633;
            10'h26f: pwm_thresh = 11'd634;
            10'h270: pwm_thresh = 11'd635;
            10'h271: pwm_thresh = 11'd636;
            10'h272: pwm_thresh = 11'd637;
            10'h273: pwm_thresh = 11'd638;
            10'h274: pwm_thresh = 11'd639;
            10'h275: pwm_thresh = 11'd640;
            10'h276: pwm_thresh = 11'd641;
            10'h277: pwm_thresh = 11'd642;
            10'h278: pwm_thresh = 11'd643;
            10'h279: pwm_thresh = 11'd644;
            10'h27a: pwm_thresh = 11'd645;
            10'h27b: pwm_thresh = 11'd646;
            10'h27c: pwm_thresh = 11'd647;
            10'h27d: pwm_thresh = 11'd648;
            10'h27e: pwm_thresh = 11'd649;
            10'h27f: pwm_thresh = 11'd650;
            10'h280: pwm_thresh = 11'd651;
            10'h281: pwm_thresh = 11'd652;
            10'h282: pwm_thresh = 11'd653;
            10'h283: pwm_thresh = 11'd654;
            10'h284: pwm_thresh = 11'd655;
            10'h285: pwm_thresh = 11'd656;
            10'h286: pwm_thresh = 11'd657;
            10'h287: pwm_thresh = 11'd659;
            10'h288: pwm_thresh = 11'd660;
            10'h289: pwm_thresh = 11'd661;
            10'h28a: pwm_thresh = 11'd662;
            10'h28b: pwm_thresh = 11'd663;
            10'h28c: pwm_thresh = 11'd664;
            10'h28d: pwm_thresh = 11'd665;
            10'h28e: pwm_thresh = 11'd666;
            10'h28f: pwm_thresh = 11'd667;
            10'h290: pwm_thresh = 11'd668;
            10'h291: pwm_thresh = 11'd669;
            10'h292: pwm_thresh = 11'd670;
            10'h293: pwm_thresh = 11'd671;
            10'h294: pwm_thresh = 11'd672;
            10'h295: pwm_thresh = 11'd673;
            10'h296: pwm_thresh = 11'd674;
            10'h297: pwm_thresh = 11'd675;
            10'h298: pwm_thresh = 11'd676;
            10'h299: pwm_thresh = 11'd677;
            10'h29a: pwm_thresh = 11'd678;
            10'h29b: pwm_thresh = 11'd679;
            10'h29c: pwm_thresh = 11'd680;
            10'h29d: pwm_thresh = 11'd681;
            10'h29e: pwm_thresh = 11'd682;
            10'h29f: pwm_thresh = 11'd683;
            10'h2a0: pwm_thresh = 11'd684;
            10'h2a1: pwm_thresh = 11'd685;
            10'h2a2: pwm_thresh = 11'd686;
            10'h2a3: pwm_thresh = 11'd687;
            10'h2a4: pwm_thresh = 11'd688;
            10'h2a5: pwm_thresh = 11'd689;
            10'h2a6: pwm_thresh = 11'd690;
            10'h2a7: pwm_thresh = 11'd691;
            10'h2a8: pwm_thresh = 11'd692;
            10'h2a9: pwm_thresh = 11'd693;
            10'h2aa: pwm_thresh = 11'd694;
            10'h2ab: pwm_thresh = 11'd695;
            10'h2ac: pwm_thresh = 11'd696;
            10'h2ad: pwm_thresh = 11'd697;
            10'h2ae: pwm_thresh = 11'd698;
            10'h2af: pwm_thresh = 11'd699;
            10'h2b0: pwm_thresh = 11'd700;
            10'h2b1: pwm_thresh = 11'd701;
            10'h2b2: pwm_thresh = 11'd702;
            10'h2b3: pwm_thresh = 11'd703;
            10'h2b4: pwm_thresh = 11'd704;
            10'h2b5: pwm_thresh = 11'd705;
            10'h2b6: pwm_thresh = 11'd706;
            10'h2b7: pwm_thresh = 11'd707;
            10'h2b8: pwm_thresh = 11'd708;
            10'h2b9: pwm_thresh = 11'd709;
            10'h2ba: pwm_thresh = 11'd710;
            10'h2bb: pwm_thresh = 11'd711;
            10'h2bc: pwm_thresh = 11'd713;
            10'h2bd: pwm_thresh = 11'd714;
            10'h2be: pwm_thresh = 11'd715;
            10'h2bf: pwm_thresh = 11'd716;
            10'h2c0: pwm_thresh = 11'd717;
            10'h2c1: pwm_thresh = 11'd718;
            10'h2c2: pwm_thresh = 11'd719;
            10'h2c3: pwm_thresh = 11'd720;
            10'h2c4: pwm_thresh = 11'd721;
            10'h2c5: pwm_thresh = 11'd722;
            10'h2c6: pwm_thresh = 11'd723;
            10'h2c7: pwm_thresh = 11'd724;
            10'h2c8: pwm_thresh = 11'd725;
            10'h2c9: pwm_thresh = 11'd726;
            10'h2ca: pwm_thresh = 11'd727;
            10'h2cb: pwm_thresh = 11'd728;
            10'h2cc: pwm_thresh = 11'd729;
            10'h2cd: pwm_thresh = 11'd730;
            10'h2ce: pwm_thresh = 11'd731;
            10'h2cf: pwm_thresh = 11'd732;
            10'h2d0: pwm_thresh = 11'd733;
            10'h2d1: pwm_thresh = 11'd734;
            10'h2d2: pwm_thresh = 11'd735;
            10'h2d3: pwm_thresh = 11'd736;
            10'h2d4: pwm_thresh = 11'd737;
            10'h2d5: pwm_thresh = 11'd738;
            10'h2d6: pwm_thresh = 11'd739;
            10'h2d7: pwm_thresh = 11'd740;
            10'h2d8: pwm_thresh = 11'd741;
            10'h2d9: pwm_thresh = 11'd742;
            10'h2da: pwm_thresh = 11'd743;
            10'h2db: pwm_thresh = 11'd744;
            10'h2dc: pwm_thresh = 11'd745;
            10'h2dd: pwm_thresh = 11'd746;
            10'h2de: pwm_thresh = 11'd747;
            10'h2df: pwm_thresh = 11'd748;
            10'h2e0: pwm_thresh = 11'd749;
            10'h2e1: pwm_thresh = 11'd750;
            10'h2e2: pwm_thresh = 11'd751;
            10'h2e3: pwm_thresh = 11'd752;
            10'h2e4: pwm_thresh = 11'd753;
            10'h2e5: pwm_thresh = 11'd754;
            10'h2e6: pwm_thresh = 11'd755;
            10'h2e7: pwm_thresh = 11'd756;
            10'h2e8: pwm_thresh = 11'd757;
            10'h2e9: pwm_thresh = 11'd758;
            10'h2ea: pwm_thresh = 11'd759;
            10'h2eb: pwm_thresh = 11'd760;
            10'h2ec: pwm_thresh = 11'd761;
            10'h2ed: pwm_thresh = 11'd762;
            10'h2ee: pwm_thresh = 11'd763;
            10'h2ef: pwm_thresh = 11'd764;
            10'h2f0: pwm_thresh = 11'd765;
            10'h2f1: pwm_thresh = 11'd766;
            10'h2f2: pwm_thresh = 11'd768;
            10'h2f3: pwm_thresh = 11'd769;
            10'h2f4: pwm_thresh = 11'd770;
            10'h2f5: pwm_thresh = 11'd771;
            10'h2f6: pwm_thresh = 11'd772;
            10'h2f7: pwm_thresh = 11'd773;
            10'h2f8: pwm_thresh = 11'd774;
            10'h2f9: pwm_thresh = 11'd775;
            10'h2fa: pwm_thresh = 11'd776;
            10'h2fb: pwm_thresh = 11'd777;
            10'h2fc: pwm_thresh = 11'd778;
            10'h2fd: pwm_thresh = 11'd779;
            10'h2fe: pwm_thresh = 11'd780;
            10'h2ff: pwm_thresh = 11'd781;
            10'h300: pwm_thresh = 11'd782;
            10'h301: pwm_thresh = 11'd783;
            10'h302: pwm_thresh = 11'd784;
            10'h303: pwm_thresh = 11'd785;
            10'h304: pwm_thresh = 11'd786;
            10'h305: pwm_thresh = 11'd787;
            10'h306: pwm_thresh = 11'd788;
            10'h307: pwm_thresh = 11'd789;
            10'h308: pwm_thresh = 11'd790;
            10'h309: pwm_thresh = 11'd791;
            10'h30a: pwm_thresh = 11'd792;
            10'h30b: pwm_thresh = 11'd793;
            10'h30c: pwm_thresh = 11'd794;
            10'h30d: pwm_thresh = 11'd795;
            10'h30e: pwm_thresh = 11'd796;
            10'h30f: pwm_thresh = 11'd797;
            10'h310: pwm_thresh = 11'd798;
            10'h311: pwm_thresh = 11'd799;
            10'h312: pwm_thresh = 11'd800;
            10'h313: pwm_thresh = 11'd801;
            10'h314: pwm_thresh = 11'd802;
            10'h315: pwm_thresh = 11'd803;
            10'h316: pwm_thresh = 11'd804;
            10'h317: pwm_thresh = 11'd805;
            10'h318: pwm_thresh = 11'd806;
            10'h319: pwm_thresh = 11'd807;
            10'h31a: pwm_thresh = 11'd808;
            10'h31b: pwm_thresh = 11'd809;
            10'h31c: pwm_thresh = 11'd810;
            10'h31d: pwm_thresh = 11'd811;
            10'h31e: pwm_thresh = 11'd812;
            10'h31f: pwm_thresh = 11'd813;
            10'h320: pwm_thresh = 11'd814;
            10'h321: pwm_thresh = 11'd815;
            10'h322: pwm_thresh = 11'd816;
            10'h323: pwm_thresh = 11'd817;
            10'h324: pwm_thresh = 11'd818;
            10'h325: pwm_thresh = 11'd819;
            10'h326: pwm_thresh = 11'd820;
            10'h327: pwm_thresh = 11'd821;
            10'h328: pwm_thresh = 11'd823;
            10'h329: pwm_thresh = 11'd824;
            10'h32a: pwm_thresh = 11'd825;
            10'h32b: pwm_thresh = 11'd826;
            10'h32c: pwm_thresh = 11'd827;
            10'h32d: pwm_thresh = 11'd828;
            10'h32e: pwm_thresh = 11'd829;
            10'h32f: pwm_thresh = 11'd830;
            10'h330: pwm_thresh = 11'd831;
            10'h331: pwm_thresh = 11'd832;
            10'h332: pwm_thresh = 11'd833;
            10'h333: pwm_thresh = 11'd834;
            10'h334: pwm_thresh = 11'd835;
            10'h335: pwm_thresh = 11'd836;
            10'h336: pwm_thresh = 11'd837;
            10'h337: pwm_thresh = 11'd838;
            10'h338: pwm_thresh = 11'd839;
            10'h339: pwm_thresh = 11'd840;
            10'h33a: pwm_thresh = 11'd841;
            10'h33b: pwm_thresh = 11'd842;
            10'h33c: pwm_thresh = 11'd843;
            10'h33d: pwm_thresh = 11'd844;
            10'h33e: pwm_thresh = 11'd845;
            10'h33f: pwm_thresh = 11'd846;
            10'h340: pwm_thresh = 11'd847;
            10'h341: pwm_thresh = 11'd848;
            10'h342: pwm_thresh = 11'd849;
            10'h343: pwm_thresh = 11'd850;
            10'h344: pwm_thresh = 11'd851;
            10'h345: pwm_thresh = 11'd852;
            10'h346: pwm_thresh = 11'd853;
            10'h347: pwm_thresh = 11'd854;
            10'h348: pwm_thresh = 11'd855;
            10'h349: pwm_thresh = 11'd856;
            10'h34a: pwm_thresh = 11'd857;
            10'h34b: pwm_thresh = 11'd858;
            10'h34c: pwm_thresh = 11'd859;
            10'h34d: pwm_thresh = 11'd860;
            10'h34e: pwm_thresh = 11'd861;
            10'h34f: pwm_thresh = 11'd862;
            10'h350: pwm_thresh = 11'd863;
            10'h351: pwm_thresh = 11'd864;
            10'h352: pwm_thresh = 11'd865;
            10'h353: pwm_thresh = 11'd866;
            10'h354: pwm_thresh = 11'd867;
            10'h355: pwm_thresh = 11'd868;
            10'h356: pwm_thresh = 11'd869;
            10'h357: pwm_thresh = 11'd870;
            10'h358: pwm_thresh = 11'd871;
            10'h359: pwm_thresh = 11'd872;
            10'h35a: pwm_thresh = 11'd873;
            10'h35b: pwm_thresh = 11'd874;
            10'h35c: pwm_thresh = 11'd875;
            10'h35d: pwm_thresh = 11'd876;
            10'h35e: pwm_thresh = 11'd878;
            10'h35f: pwm_thresh = 11'd879;
            10'h360: pwm_thresh = 11'd880;
            10'h361: pwm_thresh = 11'd881;
            10'h362: pwm_thresh = 11'd882;
            10'h363: pwm_thresh = 11'd883;
            10'h364: pwm_thresh = 11'd884;
            10'h365: pwm_thresh = 11'd885;
            10'h366: pwm_thresh = 11'd886;
            10'h367: pwm_thresh = 11'd887;
            10'h368: pwm_thresh = 11'd888;
            10'h369: pwm_thresh = 11'd889;
            10'h36a: pwm_thresh = 11'd890;
            10'h36b: pwm_thresh = 11'd891;
            10'h36c: pwm_thresh = 11'd892;
            10'h36d: pwm_thresh = 11'd893;
            10'h36e: pwm_thresh = 11'd894;
            10'h36f: pwm_thresh = 11'd895;
            10'h370: pwm_thresh = 11'd896;
            10'h371: pwm_thresh = 11'd897;
            10'h372: pwm_thresh = 11'd898;
            10'h373: pwm_thresh = 11'd899;
            10'h374: pwm_thresh = 11'd900;
            10'h375: pwm_thresh = 11'd901;
            10'h376: pwm_thresh = 11'd902;
            10'h377: pwm_thresh = 11'd903;
            10'h378: pwm_thresh = 11'd904;
            10'h379: pwm_thresh = 11'd905;
            10'h37a: pwm_thresh = 11'd906;
            10'h37b: pwm_thresh = 11'd907;
            10'h37c: pwm_thresh = 11'd908;
            10'h37d: pwm_thresh = 11'd909;
            10'h37e: pwm_thresh = 11'd910;
            10'h37f: pwm_thresh = 11'd911;
            10'h380: pwm_thresh = 11'd912;
            10'h381: pwm_thresh = 11'd913;
            10'h382: pwm_thresh = 11'd914;
            10'h383: pwm_thresh = 11'd915;
            10'h384: pwm_thresh = 11'd916;
            10'h385: pwm_thresh = 11'd917;
            10'h386: pwm_thresh = 11'd918;
            10'h387: pwm_thresh = 11'd919;
            10'h388: pwm_thresh = 11'd920;
            10'h389: pwm_thresh = 11'd921;
            10'h38a: pwm_thresh = 11'd922;
            10'h38b: pwm_thresh = 11'd923;
            10'h38c: pwm_thresh = 11'd924;
            10'h38d: pwm_thresh = 11'd925;
            10'h38e: pwm_thresh = 11'd926;
            10'h38f: pwm_thresh = 11'd927;
            10'h390: pwm_thresh = 11'd928;
            10'h391: pwm_thresh = 11'd929;
            10'h392: pwm_thresh = 11'd930;
            10'h393: pwm_thresh = 11'd931;
            10'h394: pwm_thresh = 11'd933;
            10'h395: pwm_thresh = 11'd934;
            10'h396: pwm_thresh = 11'd935;
            10'h397: pwm_thresh = 11'd936;
            10'h398: pwm_thresh = 11'd937;
            10'h399: pwm_thresh = 11'd938;
            10'h39a: pwm_thresh = 11'd939;
            10'h39b: pwm_thresh = 11'd940;
            10'h39c: pwm_thresh = 11'd941;
            10'h39d: pwm_thresh = 11'd942;
            10'h39e: pwm_thresh = 11'd943;
            10'h39f: pwm_thresh = 11'd944;
            10'h3a0: pwm_thresh = 11'd945;
            10'h3a1: pwm_thresh = 11'd946;
            10'h3a2: pwm_thresh = 11'd947;
            10'h3a3: pwm_thresh = 11'd948;
            10'h3a4: pwm_thresh = 11'd949;
            10'h3a5: pwm_thresh = 11'd950;
            10'h3a6: pwm_thresh = 11'd951;
            10'h3a7: pwm_thresh = 11'd952;
            10'h3a8: pwm_thresh = 11'd953;
            10'h3a9: pwm_thresh = 11'd954;
            10'h3aa: pwm_thresh = 11'd955;
            10'h3ab: pwm_thresh = 11'd956;
            10'h3ac: pwm_thresh = 11'd957;
            10'h3ad: pwm_thresh = 11'd958;
            10'h3ae: pwm_thresh = 11'd959;
            10'h3af: pwm_thresh = 11'd960;
            10'h3b0: pwm_thresh = 11'd961;
            10'h3b1: pwm_thresh = 11'd962;
            10'h3b2: pwm_thresh = 11'd963;
            10'h3b3: pwm_thresh = 11'd964;
            10'h3b4: pwm_thresh = 11'd965;
            10'h3b5: pwm_thresh = 11'd966;
            10'h3b6: pwm_thresh = 11'd967;
            10'h3b7: pwm_thresh = 11'd968;
            10'h3b8: pwm_thresh = 11'd969;
            10'h3b9: pwm_thresh = 11'd970;
            10'h3ba: pwm_thresh = 11'd971;
            10'h3bb: pwm_thresh = 11'd972;
            10'h3bc: pwm_thresh = 11'd973;
            10'h3bd: pwm_thresh = 11'd974;
            10'h3be: pwm_thresh = 11'd975;
            10'h3bf: pwm_thresh = 11'd976;
            10'h3c0: pwm_thresh = 11'd977;
            10'h3c1: pwm_thresh = 11'd978;
            10'h3c2: pwm_thresh = 11'd979;
            10'h3c3: pwm_thresh = 11'd980;
            10'h3c4: pwm_thresh = 11'd981;
            10'h3c5: pwm_thresh = 11'd982;
            10'h3c6: pwm_thresh = 11'd983;
            10'h3c7: pwm_thresh = 11'd984;
            10'h3c8: pwm_thresh = 11'd985;
            10'h3c9: pwm_thresh = 11'd986;
            10'h3ca: pwm_thresh = 11'd988;
            10'h3cb: pwm_thresh = 11'd989;
            10'h3cc: pwm_thresh = 11'd990;
            10'h3cd: pwm_thresh = 11'd991;
            10'h3ce: pwm_thresh = 11'd992;
            10'h3cf: pwm_thresh = 11'd993;
            10'h3d0: pwm_thresh = 11'd994;
            10'h3d1: pwm_thresh = 11'd995;
            10'h3d2: pwm_thresh = 11'd996;
            10'h3d3: pwm_thresh = 11'd997;
            10'h3d4: pwm_thresh = 11'd998;
            10'h3d5: pwm_thresh = 11'd999;
            10'h3d6: pwm_thresh = 11'd1000;
            10'h3d7: pwm_thresh = 11'd1001;
            10'h3d8: pwm_thresh = 11'd1002;
            10'h3d9: pwm_thresh = 11'd1003;
            10'h3da: pwm_thresh = 11'd1004;
            10'h3db: pwm_thresh = 11'd1005;
            10'h3dc: pwm_thresh = 11'd1006;
            10'h3dd: pwm_thresh = 11'd1007;
            10'h3de: pwm_thresh = 11'd1008;
            10'h3df: pwm_thresh = 11'd1009;
            10'h3e0: pwm_thresh = 11'd1010;
            10'h3e1: pwm_thresh = 11'd1011;
            10'h3e2: pwm_thresh = 11'd1012;
            10'h3e3: pwm_thresh = 11'd1013;
            10'h3e4: pwm_thresh = 11'd1014;
            10'h3e5: pwm_thresh = 11'd1015;
            10'h3e6: pwm_thresh = 11'd1016;
            10'h3e7: pwm_thresh = 11'd1017;
            10'h3e8: pwm_thresh = 11'd1018;
            10'h3e9: pwm_thresh = 11'd1019;
            10'h3ea: pwm_thresh = 11'd1020;
            10'h3eb: pwm_thresh = 11'd1021;
            10'h3ec: pwm_thresh = 11'd1022;
            10'h3ed: pwm_thresh = 11'd1023;
            10'h3ee: pwm_thresh = 11'd1024;
            10'h3ef: pwm_thresh = 11'd1025;
            10'h3f0: pwm_thresh = 11'd1026;
            10'h3f1: pwm_thresh = 11'd1027;
            10'h3f2: pwm_thresh = 11'd1028;
            10'h3f3: pwm_thresh = 11'd1029;
            10'h3f4: pwm_thresh = 11'd1030;
            10'h3f5: pwm_thresh = 11'd1031;
            10'h3f6: pwm_thresh = 11'd1032;
            10'h3f7: pwm_thresh = 11'd1033;
            10'h3f8: pwm_thresh = 11'd1034;
            10'h3f9: pwm_thresh = 11'd1035;
            10'h3fa: pwm_thresh = 11'd1036;
            10'h3fb: pwm_thresh = 11'd1037;
            10'h3fc: pwm_thresh = 11'd1038;
            10'h3fd: pwm_thresh = 11'd1039;
            10'h3fe: pwm_thresh = 11'd1040;
            10'h3ff: pwm_thresh = 11'd1042;
        endcase
    end

endmodule: pwm_thresh_96k
