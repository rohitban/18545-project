

module pwm_thresh_father
  (input  logic [9:0] mult_val,
   output logic [13:0] pwm_thresh);

  always_comb begin
    case(mult_val)
        10'h0: pwm_thresh = 14'd0;
        10'h1: pwm_thresh = 14'd8;
        10'h2: pwm_thresh = 14'd17;
        10'h3: pwm_thresh = 14'd26;
        10'h4: pwm_thresh = 14'd35;
        10'h5: pwm_thresh = 14'd44;
        10'h6: pwm_thresh = 14'd53;
        10'h7: pwm_thresh = 14'd62;
        10'h8: pwm_thresh = 14'd70;
        10'h9: pwm_thresh = 14'd79;
        10'ha: pwm_thresh = 14'd88;
        10'hb: pwm_thresh = 14'd97;
        10'hc: pwm_thresh = 14'd106;
        10'hd: pwm_thresh = 14'd115;
        10'he: pwm_thresh = 14'd124;
        10'hf: pwm_thresh = 14'd132;
        10'h10: pwm_thresh = 14'd141;
        10'h11: pwm_thresh = 14'd150;
        10'h12: pwm_thresh = 14'd159;
        10'h13: pwm_thresh = 14'd168;
        10'h14: pwm_thresh = 14'd177;
        10'h15: pwm_thresh = 14'd186;
        10'h16: pwm_thresh = 14'd195;
        10'h17: pwm_thresh = 14'd203;
        10'h18: pwm_thresh = 14'd212;
        10'h19: pwm_thresh = 14'd221;
        10'h1a: pwm_thresh = 14'd230;
        10'h1b: pwm_thresh = 14'd239;
        10'h1c: pwm_thresh = 14'd248;
        10'h1d: pwm_thresh = 14'd257;
        10'h1e: pwm_thresh = 14'd265;
        10'h1f: pwm_thresh = 14'd274;
        10'h20: pwm_thresh = 14'd283;
        10'h21: pwm_thresh = 14'd292;
        10'h22: pwm_thresh = 14'd301;
        10'h23: pwm_thresh = 14'd310;
        10'h24: pwm_thresh = 14'd319;
        10'h25: pwm_thresh = 14'd328;
        10'h26: pwm_thresh = 14'd336;
        10'h27: pwm_thresh = 14'd345;
        10'h28: pwm_thresh = 14'd354;
        10'h29: pwm_thresh = 14'd363;
        10'h2a: pwm_thresh = 14'd372;
        10'h2b: pwm_thresh = 14'd381;
        10'h2c: pwm_thresh = 14'd390;
        10'h2d: pwm_thresh = 14'd398;
        10'h2e: pwm_thresh = 14'd407;
        10'h2f: pwm_thresh = 14'd416;
        10'h30: pwm_thresh = 14'd425;
        10'h31: pwm_thresh = 14'd434;
        10'h32: pwm_thresh = 14'd443;
        10'h33: pwm_thresh = 14'd452;
        10'h34: pwm_thresh = 14'd461;
        10'h35: pwm_thresh = 14'd469;
        10'h36: pwm_thresh = 14'd478;
        10'h37: pwm_thresh = 14'd487;
        10'h38: pwm_thresh = 14'd496;
        10'h39: pwm_thresh = 14'd505;
        10'h3a: pwm_thresh = 14'd514;
        10'h3b: pwm_thresh = 14'd523;
        10'h3c: pwm_thresh = 14'd531;
        10'h3d: pwm_thresh = 14'd540;
        10'h3e: pwm_thresh = 14'd549;
        10'h3f: pwm_thresh = 14'd558;
        10'h40: pwm_thresh = 14'd567;
        10'h41: pwm_thresh = 14'd576;
        10'h42: pwm_thresh = 14'd585;
        10'h43: pwm_thresh = 14'd594;
        10'h44: pwm_thresh = 14'd602;
        10'h45: pwm_thresh = 14'd611;
        10'h46: pwm_thresh = 14'd620;
        10'h47: pwm_thresh = 14'd629;
        10'h48: pwm_thresh = 14'd638;
        10'h49: pwm_thresh = 14'd647;
        10'h4a: pwm_thresh = 14'd656;
        10'h4b: pwm_thresh = 14'd664;
        10'h4c: pwm_thresh = 14'd673;
        10'h4d: pwm_thresh = 14'd682;
        10'h4e: pwm_thresh = 14'd691;
        10'h4f: pwm_thresh = 14'd700;
        10'h50: pwm_thresh = 14'd709;
        10'h51: pwm_thresh = 14'd718;
        10'h52: pwm_thresh = 14'd727;
        10'h53: pwm_thresh = 14'd735;
        10'h54: pwm_thresh = 14'd744;
        10'h55: pwm_thresh = 14'd753;
        10'h56: pwm_thresh = 14'd762;
        10'h57: pwm_thresh = 14'd771;
        10'h58: pwm_thresh = 14'd780;
        10'h59: pwm_thresh = 14'd789;
        10'h5a: pwm_thresh = 14'd797;
        10'h5b: pwm_thresh = 14'd806;
        10'h5c: pwm_thresh = 14'd815;
        10'h5d: pwm_thresh = 14'd824;
        10'h5e: pwm_thresh = 14'd833;
        10'h5f: pwm_thresh = 14'd842;
        10'h60: pwm_thresh = 14'd851;
        10'h61: pwm_thresh = 14'd860;
        10'h62: pwm_thresh = 14'd868;
        10'h63: pwm_thresh = 14'd877;
        10'h64: pwm_thresh = 14'd886;
        10'h65: pwm_thresh = 14'd895;
        10'h66: pwm_thresh = 14'd904;
        10'h67: pwm_thresh = 14'd913;
        10'h68: pwm_thresh = 14'd922;
        10'h69: pwm_thresh = 14'd930;
        10'h6a: pwm_thresh = 14'd939;
        10'h6b: pwm_thresh = 14'd948;
        10'h6c: pwm_thresh = 14'd957;
        10'h6d: pwm_thresh = 14'd966;
        10'h6e: pwm_thresh = 14'd975;
        10'h6f: pwm_thresh = 14'd984;
        10'h70: pwm_thresh = 14'd993;
        10'h71: pwm_thresh = 14'd1001;
        10'h72: pwm_thresh = 14'd1010;
        10'h73: pwm_thresh = 14'd1019;
        10'h74: pwm_thresh = 14'd1028;
        10'h75: pwm_thresh = 14'd1037;
        10'h76: pwm_thresh = 14'd1046;
        10'h77: pwm_thresh = 14'd1055;
        10'h78: pwm_thresh = 14'd1063;
        10'h79: pwm_thresh = 14'd1072;
        10'h7a: pwm_thresh = 14'd1081;
        10'h7b: pwm_thresh = 14'd1090;
        10'h7c: pwm_thresh = 14'd1099;
        10'h7d: pwm_thresh = 14'd1108;
        10'h7e: pwm_thresh = 14'd1117;
        10'h7f: pwm_thresh = 14'd1125;
        10'h80: pwm_thresh = 14'd1134;
        10'h81: pwm_thresh = 14'd1143;
        10'h82: pwm_thresh = 14'd1152;
        10'h83: pwm_thresh = 14'd1161;
        10'h84: pwm_thresh = 14'd1170;
        10'h85: pwm_thresh = 14'd1179;
        10'h86: pwm_thresh = 14'd1188;
        10'h87: pwm_thresh = 14'd1196;
        10'h88: pwm_thresh = 14'd1205;
        10'h89: pwm_thresh = 14'd1214;
        10'h8a: pwm_thresh = 14'd1223;
        10'h8b: pwm_thresh = 14'd1232;
        10'h8c: pwm_thresh = 14'd1241;
        10'h8d: pwm_thresh = 14'd1250;
        10'h8e: pwm_thresh = 14'd1258;
        10'h8f: pwm_thresh = 14'd1267;
        10'h90: pwm_thresh = 14'd1276;
        10'h91: pwm_thresh = 14'd1285;
        10'h92: pwm_thresh = 14'd1294;
        10'h93: pwm_thresh = 14'd1303;
        10'h94: pwm_thresh = 14'd1312;
        10'h95: pwm_thresh = 14'd1321;
        10'h96: pwm_thresh = 14'd1329;
        10'h97: pwm_thresh = 14'd1338;
        10'h98: pwm_thresh = 14'd1347;
        10'h99: pwm_thresh = 14'd1356;
        10'h9a: pwm_thresh = 14'd1365;
        10'h9b: pwm_thresh = 14'd1374;
        10'h9c: pwm_thresh = 14'd1383;
        10'h9d: pwm_thresh = 14'd1391;
        10'h9e: pwm_thresh = 14'd1400;
        10'h9f: pwm_thresh = 14'd1409;
        10'ha0: pwm_thresh = 14'd1418;
        10'ha1: pwm_thresh = 14'd1427;
        10'ha2: pwm_thresh = 14'd1436;
        10'ha3: pwm_thresh = 14'd1445;
        10'ha4: pwm_thresh = 14'd1454;
        10'ha5: pwm_thresh = 14'd1462;
        10'ha6: pwm_thresh = 14'd1471;
        10'ha7: pwm_thresh = 14'd1480;
        10'ha8: pwm_thresh = 14'd1489;
        10'ha9: pwm_thresh = 14'd1498;
        10'haa: pwm_thresh = 14'd1507;
        10'hab: pwm_thresh = 14'd1516;
        10'hac: pwm_thresh = 14'd1524;
        10'had: pwm_thresh = 14'd1533;
        10'hae: pwm_thresh = 14'd1542;
        10'haf: pwm_thresh = 14'd1551;
        10'hb0: pwm_thresh = 14'd1560;
        10'hb1: pwm_thresh = 14'd1569;
        10'hb2: pwm_thresh = 14'd1578;
        10'hb3: pwm_thresh = 14'd1587;
        10'hb4: pwm_thresh = 14'd1595;
        10'hb5: pwm_thresh = 14'd1604;
        10'hb6: pwm_thresh = 14'd1613;
        10'hb7: pwm_thresh = 14'd1622;
        10'hb8: pwm_thresh = 14'd1631;
        10'hb9: pwm_thresh = 14'd1640;
        10'hba: pwm_thresh = 14'd1649;
        10'hbb: pwm_thresh = 14'd1657;
        10'hbc: pwm_thresh = 14'd1666;
        10'hbd: pwm_thresh = 14'd1675;
        10'hbe: pwm_thresh = 14'd1684;
        10'hbf: pwm_thresh = 14'd1693;
        10'hc0: pwm_thresh = 14'd1702;
        10'hc1: pwm_thresh = 14'd1711;
        10'hc2: pwm_thresh = 14'd1720;
        10'hc3: pwm_thresh = 14'd1728;
        10'hc4: pwm_thresh = 14'd1737;
        10'hc5: pwm_thresh = 14'd1746;
        10'hc6: pwm_thresh = 14'd1755;
        10'hc7: pwm_thresh = 14'd1764;
        10'hc8: pwm_thresh = 14'd1773;
        10'hc9: pwm_thresh = 14'd1782;
        10'hca: pwm_thresh = 14'd1790;
        10'hcb: pwm_thresh = 14'd1799;
        10'hcc: pwm_thresh = 14'd1808;
        10'hcd: pwm_thresh = 14'd1817;
        10'hce: pwm_thresh = 14'd1826;
        10'hcf: pwm_thresh = 14'd1835;
        10'hd0: pwm_thresh = 14'd1844;
        10'hd1: pwm_thresh = 14'd1853;
        10'hd2: pwm_thresh = 14'd1861;
        10'hd3: pwm_thresh = 14'd1870;
        10'hd4: pwm_thresh = 14'd1879;
        10'hd5: pwm_thresh = 14'd1888;
        10'hd6: pwm_thresh = 14'd1897;
        10'hd7: pwm_thresh = 14'd1906;
        10'hd8: pwm_thresh = 14'd1915;
        10'hd9: pwm_thresh = 14'd1923;
        10'hda: pwm_thresh = 14'd1932;
        10'hdb: pwm_thresh = 14'd1941;
        10'hdc: pwm_thresh = 14'd1950;
        10'hdd: pwm_thresh = 14'd1959;
        10'hde: pwm_thresh = 14'd1968;
        10'hdf: pwm_thresh = 14'd1977;
        10'he0: pwm_thresh = 14'd1986;
        10'he1: pwm_thresh = 14'd1994;
        10'he2: pwm_thresh = 14'd2003;
        10'he3: pwm_thresh = 14'd2012;
        10'he4: pwm_thresh = 14'd2021;
        10'he5: pwm_thresh = 14'd2030;
        10'he6: pwm_thresh = 14'd2039;
        10'he7: pwm_thresh = 14'd2048;
        10'he8: pwm_thresh = 14'd2056;
        10'he9: pwm_thresh = 14'd2065;
        10'hea: pwm_thresh = 14'd2074;
        10'heb: pwm_thresh = 14'd2083;
        10'hec: pwm_thresh = 14'd2092;
        10'hed: pwm_thresh = 14'd2101;
        10'hee: pwm_thresh = 14'd2110;
        10'hef: pwm_thresh = 14'd2118;
        10'hf0: pwm_thresh = 14'd2127;
        10'hf1: pwm_thresh = 14'd2136;
        10'hf2: pwm_thresh = 14'd2145;
        10'hf3: pwm_thresh = 14'd2154;
        10'hf4: pwm_thresh = 14'd2163;
        10'hf5: pwm_thresh = 14'd2172;
        10'hf6: pwm_thresh = 14'd2181;
        10'hf7: pwm_thresh = 14'd2189;
        10'hf8: pwm_thresh = 14'd2198;
        10'hf9: pwm_thresh = 14'd2207;
        10'hfa: pwm_thresh = 14'd2216;
        10'hfb: pwm_thresh = 14'd2225;
        10'hfc: pwm_thresh = 14'd2234;
        10'hfd: pwm_thresh = 14'd2243;
        10'hfe: pwm_thresh = 14'd2251;
        10'hff: pwm_thresh = 14'd2260;
        10'h100: pwm_thresh = 14'd2269;
        10'h101: pwm_thresh = 14'd2278;
        10'h102: pwm_thresh = 14'd2287;
        10'h103: pwm_thresh = 14'd2296;
        10'h104: pwm_thresh = 14'd2305;
        10'h105: pwm_thresh = 14'd2314;
        10'h106: pwm_thresh = 14'd2322;
        10'h107: pwm_thresh = 14'd2331;
        10'h108: pwm_thresh = 14'd2340;
        10'h109: pwm_thresh = 14'd2349;
        10'h10a: pwm_thresh = 14'd2358;
        10'h10b: pwm_thresh = 14'd2367;
        10'h10c: pwm_thresh = 14'd2376;
        10'h10d: pwm_thresh = 14'd2384;
        10'h10e: pwm_thresh = 14'd2393;
        10'h10f: pwm_thresh = 14'd2402;
        10'h110: pwm_thresh = 14'd2411;
        10'h111: pwm_thresh = 14'd2420;
        10'h112: pwm_thresh = 14'd2429;
        10'h113: pwm_thresh = 14'd2438;
        10'h114: pwm_thresh = 14'd2447;
        10'h115: pwm_thresh = 14'd2455;
        10'h116: pwm_thresh = 14'd2464;
        10'h117: pwm_thresh = 14'd2473;
        10'h118: pwm_thresh = 14'd2482;
        10'h119: pwm_thresh = 14'd2491;
        10'h11a: pwm_thresh = 14'd2500;
        10'h11b: pwm_thresh = 14'd2509;
        10'h11c: pwm_thresh = 14'd2517;
        10'h11d: pwm_thresh = 14'd2526;
        10'h11e: pwm_thresh = 14'd2535;
        10'h11f: pwm_thresh = 14'd2544;
        10'h120: pwm_thresh = 14'd2553;
        10'h121: pwm_thresh = 14'd2562;
        10'h122: pwm_thresh = 14'd2571;
        10'h123: pwm_thresh = 14'd2580;
        10'h124: pwm_thresh = 14'd2588;
        10'h125: pwm_thresh = 14'd2597;
        10'h126: pwm_thresh = 14'd2606;
        10'h127: pwm_thresh = 14'd2615;
        10'h128: pwm_thresh = 14'd2624;
        10'h129: pwm_thresh = 14'd2633;
        10'h12a: pwm_thresh = 14'd2642;
        10'h12b: pwm_thresh = 14'd2650;
        10'h12c: pwm_thresh = 14'd2659;
        10'h12d: pwm_thresh = 14'd2668;
        10'h12e: pwm_thresh = 14'd2677;
        10'h12f: pwm_thresh = 14'd2686;
        10'h130: pwm_thresh = 14'd2695;
        10'h131: pwm_thresh = 14'd2704;
        10'h132: pwm_thresh = 14'd2713;
        10'h133: pwm_thresh = 14'd2721;
        10'h134: pwm_thresh = 14'd2730;
        10'h135: pwm_thresh = 14'd2739;
        10'h136: pwm_thresh = 14'd2748;
        10'h137: pwm_thresh = 14'd2757;
        10'h138: pwm_thresh = 14'd2766;
        10'h139: pwm_thresh = 14'd2775;
        10'h13a: pwm_thresh = 14'd2783;
        10'h13b: pwm_thresh = 14'd2792;
        10'h13c: pwm_thresh = 14'd2801;
        10'h13d: pwm_thresh = 14'd2810;
        10'h13e: pwm_thresh = 14'd2819;
        10'h13f: pwm_thresh = 14'd2828;
        10'h140: pwm_thresh = 14'd2837;
        10'h141: pwm_thresh = 14'd2846;
        10'h142: pwm_thresh = 14'd2854;
        10'h143: pwm_thresh = 14'd2863;
        10'h144: pwm_thresh = 14'd2872;
        10'h145: pwm_thresh = 14'd2881;
        10'h146: pwm_thresh = 14'd2890;
        10'h147: pwm_thresh = 14'd2899;
        10'h148: pwm_thresh = 14'd2908;
        10'h149: pwm_thresh = 14'd2916;
        10'h14a: pwm_thresh = 14'd2925;
        10'h14b: pwm_thresh = 14'd2934;
        10'h14c: pwm_thresh = 14'd2943;
        10'h14d: pwm_thresh = 14'd2952;
        10'h14e: pwm_thresh = 14'd2961;
        10'h14f: pwm_thresh = 14'd2970;
        10'h150: pwm_thresh = 14'd2979;
        10'h151: pwm_thresh = 14'd2987;
        10'h152: pwm_thresh = 14'd2996;
        10'h153: pwm_thresh = 14'd3005;
        10'h154: pwm_thresh = 14'd3014;
        10'h155: pwm_thresh = 14'd3023;
        10'h156: pwm_thresh = 14'd3032;
        10'h157: pwm_thresh = 14'd3041;
        10'h158: pwm_thresh = 14'd3049;
        10'h159: pwm_thresh = 14'd3058;
        10'h15a: pwm_thresh = 14'd3067;
        10'h15b: pwm_thresh = 14'd3076;
        10'h15c: pwm_thresh = 14'd3085;
        10'h15d: pwm_thresh = 14'd3094;
        10'h15e: pwm_thresh = 14'd3103;
        10'h15f: pwm_thresh = 14'd3111;
        10'h160: pwm_thresh = 14'd3120;
        10'h161: pwm_thresh = 14'd3129;
        10'h162: pwm_thresh = 14'd3138;
        10'h163: pwm_thresh = 14'd3147;
        10'h164: pwm_thresh = 14'd3156;
        10'h165: pwm_thresh = 14'd3165;
        10'h166: pwm_thresh = 14'd3174;
        10'h167: pwm_thresh = 14'd3182;
        10'h168: pwm_thresh = 14'd3191;
        10'h169: pwm_thresh = 14'd3200;
        10'h16a: pwm_thresh = 14'd3209;
        10'h16b: pwm_thresh = 14'd3218;
        10'h16c: pwm_thresh = 14'd3227;
        10'h16d: pwm_thresh = 14'd3236;
        10'h16e: pwm_thresh = 14'd3244;
        10'h16f: pwm_thresh = 14'd3253;
        10'h170: pwm_thresh = 14'd3262;
        10'h171: pwm_thresh = 14'd3271;
        10'h172: pwm_thresh = 14'd3280;
        10'h173: pwm_thresh = 14'd3289;
        10'h174: pwm_thresh = 14'd3298;
        10'h175: pwm_thresh = 14'd3307;
        10'h176: pwm_thresh = 14'd3315;
        10'h177: pwm_thresh = 14'd3324;
        10'h178: pwm_thresh = 14'd3333;
        10'h179: pwm_thresh = 14'd3342;
        10'h17a: pwm_thresh = 14'd3351;
        10'h17b: pwm_thresh = 14'd3360;
        10'h17c: pwm_thresh = 14'd3369;
        10'h17d: pwm_thresh = 14'd3377;
        10'h17e: pwm_thresh = 14'd3386;
        10'h17f: pwm_thresh = 14'd3395;
        10'h180: pwm_thresh = 14'd3404;
        10'h181: pwm_thresh = 14'd3413;
        10'h182: pwm_thresh = 14'd3422;
        10'h183: pwm_thresh = 14'd3431;
        10'h184: pwm_thresh = 14'd3440;
        10'h185: pwm_thresh = 14'd3448;
        10'h186: pwm_thresh = 14'd3457;
        10'h187: pwm_thresh = 14'd3466;
        10'h188: pwm_thresh = 14'd3475;
        10'h189: pwm_thresh = 14'd3484;
        10'h18a: pwm_thresh = 14'd3493;
        10'h18b: pwm_thresh = 14'd3502;
        10'h18c: pwm_thresh = 14'd3510;
        10'h18d: pwm_thresh = 14'd3519;
        10'h18e: pwm_thresh = 14'd3528;
        10'h18f: pwm_thresh = 14'd3537;
        10'h190: pwm_thresh = 14'd3546;
        10'h191: pwm_thresh = 14'd3555;
        10'h192: pwm_thresh = 14'd3564;
        10'h193: pwm_thresh = 14'd3573;
        10'h194: pwm_thresh = 14'd3581;
        10'h195: pwm_thresh = 14'd3590;
        10'h196: pwm_thresh = 14'd3599;
        10'h197: pwm_thresh = 14'd3608;
        10'h198: pwm_thresh = 14'd3617;
        10'h199: pwm_thresh = 14'd3626;
        10'h19a: pwm_thresh = 14'd3635;
        10'h19b: pwm_thresh = 14'd3643;
        10'h19c: pwm_thresh = 14'd3652;
        10'h19d: pwm_thresh = 14'd3661;
        10'h19e: pwm_thresh = 14'd3670;
        10'h19f: pwm_thresh = 14'd3679;
        10'h1a0: pwm_thresh = 14'd3688;
        10'h1a1: pwm_thresh = 14'd3697;
        10'h1a2: pwm_thresh = 14'd3706;
        10'h1a3: pwm_thresh = 14'd3714;
        10'h1a4: pwm_thresh = 14'd3723;
        10'h1a5: pwm_thresh = 14'd3732;
        10'h1a6: pwm_thresh = 14'd3741;
        10'h1a7: pwm_thresh = 14'd3750;
        10'h1a8: pwm_thresh = 14'd3759;
        10'h1a9: pwm_thresh = 14'd3768;
        10'h1aa: pwm_thresh = 14'd3776;
        10'h1ab: pwm_thresh = 14'd3785;
        10'h1ac: pwm_thresh = 14'd3794;
        10'h1ad: pwm_thresh = 14'd3803;
        10'h1ae: pwm_thresh = 14'd3812;
        10'h1af: pwm_thresh = 14'd3821;
        10'h1b0: pwm_thresh = 14'd3830;
        10'h1b1: pwm_thresh = 14'd3839;
        10'h1b2: pwm_thresh = 14'd3847;
        10'h1b3: pwm_thresh = 14'd3856;
        10'h1b4: pwm_thresh = 14'd3865;
        10'h1b5: pwm_thresh = 14'd3874;
        10'h1b6: pwm_thresh = 14'd3883;
        10'h1b7: pwm_thresh = 14'd3892;
        10'h1b8: pwm_thresh = 14'd3901;
        10'h1b9: pwm_thresh = 14'd3909;
        10'h1ba: pwm_thresh = 14'd3918;
        10'h1bb: pwm_thresh = 14'd3927;
        10'h1bc: pwm_thresh = 14'd3936;
        10'h1bd: pwm_thresh = 14'd3945;
        10'h1be: pwm_thresh = 14'd3954;
        10'h1bf: pwm_thresh = 14'd3963;
        10'h1c0: pwm_thresh = 14'd3972;
        10'h1c1: pwm_thresh = 14'd3980;
        10'h1c2: pwm_thresh = 14'd3989;
        10'h1c3: pwm_thresh = 14'd3998;
        10'h1c4: pwm_thresh = 14'd4007;
        10'h1c5: pwm_thresh = 14'd4016;
        10'h1c6: pwm_thresh = 14'd4025;
        10'h1c7: pwm_thresh = 14'd4034;
        10'h1c8: pwm_thresh = 14'd4042;
        10'h1c9: pwm_thresh = 14'd4051;
        10'h1ca: pwm_thresh = 14'd4060;
        10'h1cb: pwm_thresh = 14'd4069;
        10'h1cc: pwm_thresh = 14'd4078;
        10'h1cd: pwm_thresh = 14'd4087;
        10'h1ce: pwm_thresh = 14'd4096;
        10'h1cf: pwm_thresh = 14'd4104;
        10'h1d0: pwm_thresh = 14'd4113;
        10'h1d1: pwm_thresh = 14'd4122;
        10'h1d2: pwm_thresh = 14'd4131;
        10'h1d3: pwm_thresh = 14'd4140;
        10'h1d4: pwm_thresh = 14'd4149;
        10'h1d5: pwm_thresh = 14'd4158;
        10'h1d6: pwm_thresh = 14'd4167;
        10'h1d7: pwm_thresh = 14'd4175;
        10'h1d8: pwm_thresh = 14'd4184;
        10'h1d9: pwm_thresh = 14'd4193;
        10'h1da: pwm_thresh = 14'd4202;
        10'h1db: pwm_thresh = 14'd4211;
        10'h1dc: pwm_thresh = 14'd4220;
        10'h1dd: pwm_thresh = 14'd4229;
        10'h1de: pwm_thresh = 14'd4237;
        10'h1df: pwm_thresh = 14'd4246;
        10'h1e0: pwm_thresh = 14'd4255;
        10'h1e1: pwm_thresh = 14'd4264;
        10'h1e2: pwm_thresh = 14'd4273;
        10'h1e3: pwm_thresh = 14'd4282;
        10'h1e4: pwm_thresh = 14'd4291;
        10'h1e5: pwm_thresh = 14'd4300;
        10'h1e6: pwm_thresh = 14'd4308;
        10'h1e7: pwm_thresh = 14'd4317;
        10'h1e8: pwm_thresh = 14'd4326;
        10'h1e9: pwm_thresh = 14'd4335;
        10'h1ea: pwm_thresh = 14'd4344;
        10'h1eb: pwm_thresh = 14'd4353;
        10'h1ec: pwm_thresh = 14'd4362;
        10'h1ed: pwm_thresh = 14'd4370;
        10'h1ee: pwm_thresh = 14'd4379;
        10'h1ef: pwm_thresh = 14'd4388;
        10'h1f0: pwm_thresh = 14'd4397;
        10'h1f1: pwm_thresh = 14'd4406;
        10'h1f2: pwm_thresh = 14'd4415;
        10'h1f3: pwm_thresh = 14'd4424;
        10'h1f4: pwm_thresh = 14'd4433;
        10'h1f5: pwm_thresh = 14'd4441;
        10'h1f6: pwm_thresh = 14'd4450;
        10'h1f7: pwm_thresh = 14'd4459;
        10'h1f8: pwm_thresh = 14'd4468;
        10'h1f9: pwm_thresh = 14'd4477;
        10'h1fa: pwm_thresh = 14'd4486;
        10'h1fb: pwm_thresh = 14'd4495;
        10'h1fc: pwm_thresh = 14'd4503;
        10'h1fd: pwm_thresh = 14'd4512;
        10'h1fe: pwm_thresh = 14'd4521;
        10'h1ff: pwm_thresh = 14'd4530;
        10'h200: pwm_thresh = 14'd4539;
        10'h201: pwm_thresh = 14'd4548;
        10'h202: pwm_thresh = 14'd4557;
        10'h203: pwm_thresh = 14'd4566;
        10'h204: pwm_thresh = 14'd4574;
        10'h205: pwm_thresh = 14'd4583;
        10'h206: pwm_thresh = 14'd4592;
        10'h207: pwm_thresh = 14'd4601;
        10'h208: pwm_thresh = 14'd4610;
        10'h209: pwm_thresh = 14'd4619;
        10'h20a: pwm_thresh = 14'd4628;
        10'h20b: pwm_thresh = 14'd4636;
        10'h20c: pwm_thresh = 14'd4645;
        10'h20d: pwm_thresh = 14'd4654;
        10'h20e: pwm_thresh = 14'd4663;
        10'h20f: pwm_thresh = 14'd4672;
        10'h210: pwm_thresh = 14'd4681;
        10'h211: pwm_thresh = 14'd4690;
        10'h212: pwm_thresh = 14'd4699;
        10'h213: pwm_thresh = 14'd4707;
        10'h214: pwm_thresh = 14'd4716;
        10'h215: pwm_thresh = 14'd4725;
        10'h216: pwm_thresh = 14'd4734;
        10'h217: pwm_thresh = 14'd4743;
        10'h218: pwm_thresh = 14'd4752;
        10'h219: pwm_thresh = 14'd4761;
        10'h21a: pwm_thresh = 14'd4769;
        10'h21b: pwm_thresh = 14'd4778;
        10'h21c: pwm_thresh = 14'd4787;
        10'h21d: pwm_thresh = 14'd4796;
        10'h21e: pwm_thresh = 14'd4805;
        10'h21f: pwm_thresh = 14'd4814;
        10'h220: pwm_thresh = 14'd4823;
        10'h221: pwm_thresh = 14'd4832;
        10'h222: pwm_thresh = 14'd4840;
        10'h223: pwm_thresh = 14'd4849;
        10'h224: pwm_thresh = 14'd4858;
        10'h225: pwm_thresh = 14'd4867;
        10'h226: pwm_thresh = 14'd4876;
        10'h227: pwm_thresh = 14'd4885;
        10'h228: pwm_thresh = 14'd4894;
        10'h229: pwm_thresh = 14'd4902;
        10'h22a: pwm_thresh = 14'd4911;
        10'h22b: pwm_thresh = 14'd4920;
        10'h22c: pwm_thresh = 14'd4929;
        10'h22d: pwm_thresh = 14'd4938;
        10'h22e: pwm_thresh = 14'd4947;
        10'h22f: pwm_thresh = 14'd4956;
        10'h230: pwm_thresh = 14'd4965;
        10'h231: pwm_thresh = 14'd4973;
        10'h232: pwm_thresh = 14'd4982;
        10'h233: pwm_thresh = 14'd4991;
        10'h234: pwm_thresh = 14'd5000;
        10'h235: pwm_thresh = 14'd5009;
        10'h236: pwm_thresh = 14'd5018;
        10'h237: pwm_thresh = 14'd5027;
        10'h238: pwm_thresh = 14'd5035;
        10'h239: pwm_thresh = 14'd5044;
        10'h23a: pwm_thresh = 14'd5053;
        10'h23b: pwm_thresh = 14'd5062;
        10'h23c: pwm_thresh = 14'd5071;
        10'h23d: pwm_thresh = 14'd5080;
        10'h23e: pwm_thresh = 14'd5089;
        10'h23f: pwm_thresh = 14'd5097;
        10'h240: pwm_thresh = 14'd5106;
        10'h241: pwm_thresh = 14'd5115;
        10'h242: pwm_thresh = 14'd5124;
        10'h243: pwm_thresh = 14'd5133;
        10'h244: pwm_thresh = 14'd5142;
        10'h245: pwm_thresh = 14'd5151;
        10'h246: pwm_thresh = 14'd5160;
        10'h247: pwm_thresh = 14'd5168;
        10'h248: pwm_thresh = 14'd5177;
        10'h249: pwm_thresh = 14'd5186;
        10'h24a: pwm_thresh = 14'd5195;
        10'h24b: pwm_thresh = 14'd5204;
        10'h24c: pwm_thresh = 14'd5213;
        10'h24d: pwm_thresh = 14'd5222;
        10'h24e: pwm_thresh = 14'd5230;
        10'h24f: pwm_thresh = 14'd5239;
        10'h250: pwm_thresh = 14'd5248;
        10'h251: pwm_thresh = 14'd5257;
        10'h252: pwm_thresh = 14'd5266;
        10'h253: pwm_thresh = 14'd5275;
        10'h254: pwm_thresh = 14'd5284;
        10'h255: pwm_thresh = 14'd5293;
        10'h256: pwm_thresh = 14'd5301;
        10'h257: pwm_thresh = 14'd5310;
        10'h258: pwm_thresh = 14'd5319;
        10'h259: pwm_thresh = 14'd5328;
        10'h25a: pwm_thresh = 14'd5337;
        10'h25b: pwm_thresh = 14'd5346;
        10'h25c: pwm_thresh = 14'd5355;
        10'h25d: pwm_thresh = 14'd5363;
        10'h25e: pwm_thresh = 14'd5372;
        10'h25f: pwm_thresh = 14'd5381;
        10'h260: pwm_thresh = 14'd5390;
        10'h261: pwm_thresh = 14'd5399;
        10'h262: pwm_thresh = 14'd5408;
        10'h263: pwm_thresh = 14'd5417;
        10'h264: pwm_thresh = 14'd5426;
        10'h265: pwm_thresh = 14'd5434;
        10'h266: pwm_thresh = 14'd5443;
        10'h267: pwm_thresh = 14'd5452;
        10'h268: pwm_thresh = 14'd5461;
        10'h269: pwm_thresh = 14'd5470;
        10'h26a: pwm_thresh = 14'd5479;
        10'h26b: pwm_thresh = 14'd5488;
        10'h26c: pwm_thresh = 14'd5496;
        10'h26d: pwm_thresh = 14'd5505;
        10'h26e: pwm_thresh = 14'd5514;
        10'h26f: pwm_thresh = 14'd5523;
        10'h270: pwm_thresh = 14'd5532;
        10'h271: pwm_thresh = 14'd5541;
        10'h272: pwm_thresh = 14'd5550;
        10'h273: pwm_thresh = 14'd5559;
        10'h274: pwm_thresh = 14'd5567;
        10'h275: pwm_thresh = 14'd5576;
        10'h276: pwm_thresh = 14'd5585;
        10'h277: pwm_thresh = 14'd5594;
        10'h278: pwm_thresh = 14'd5603;
        10'h279: pwm_thresh = 14'd5612;
        10'h27a: pwm_thresh = 14'd5621;
        10'h27b: pwm_thresh = 14'd5629;
        10'h27c: pwm_thresh = 14'd5638;
        10'h27d: pwm_thresh = 14'd5647;
        10'h27e: pwm_thresh = 14'd5656;
        10'h27f: pwm_thresh = 14'd5665;
        10'h280: pwm_thresh = 14'd5674;
        10'h281: pwm_thresh = 14'd5683;
        10'h282: pwm_thresh = 14'd5692;
        10'h283: pwm_thresh = 14'd5700;
        10'h284: pwm_thresh = 14'd5709;
        10'h285: pwm_thresh = 14'd5718;
        10'h286: pwm_thresh = 14'd5727;
        10'h287: pwm_thresh = 14'd5736;
        10'h288: pwm_thresh = 14'd5745;
        10'h289: pwm_thresh = 14'd5754;
        10'h28a: pwm_thresh = 14'd5762;
        10'h28b: pwm_thresh = 14'd5771;
        10'h28c: pwm_thresh = 14'd5780;
        10'h28d: pwm_thresh = 14'd5789;
        10'h28e: pwm_thresh = 14'd5798;
        10'h28f: pwm_thresh = 14'd5807;
        10'h290: pwm_thresh = 14'd5816;
        10'h291: pwm_thresh = 14'd5825;
        10'h292: pwm_thresh = 14'd5833;
        10'h293: pwm_thresh = 14'd5842;
        10'h294: pwm_thresh = 14'd5851;
        10'h295: pwm_thresh = 14'd5860;
        10'h296: pwm_thresh = 14'd5869;
        10'h297: pwm_thresh = 14'd5878;
        10'h298: pwm_thresh = 14'd5887;
        10'h299: pwm_thresh = 14'd5895;
        10'h29a: pwm_thresh = 14'd5904;
        10'h29b: pwm_thresh = 14'd5913;
        10'h29c: pwm_thresh = 14'd5922;
        10'h29d: pwm_thresh = 14'd5931;
        10'h29e: pwm_thresh = 14'd5940;
        10'h29f: pwm_thresh = 14'd5949;
        10'h2a0: pwm_thresh = 14'd5958;
        10'h2a1: pwm_thresh = 14'd5966;
        10'h2a2: pwm_thresh = 14'd5975;
        10'h2a3: pwm_thresh = 14'd5984;
        10'h2a4: pwm_thresh = 14'd5993;
        10'h2a5: pwm_thresh = 14'd6002;
        10'h2a6: pwm_thresh = 14'd6011;
        10'h2a7: pwm_thresh = 14'd6020;
        10'h2a8: pwm_thresh = 14'd6028;
        10'h2a9: pwm_thresh = 14'd6037;
        10'h2aa: pwm_thresh = 14'd6046;
        10'h2ab: pwm_thresh = 14'd6055;
        10'h2ac: pwm_thresh = 14'd6064;
        10'h2ad: pwm_thresh = 14'd6073;
        10'h2ae: pwm_thresh = 14'd6082;
        10'h2af: pwm_thresh = 14'd6090;
        10'h2b0: pwm_thresh = 14'd6099;
        10'h2b1: pwm_thresh = 14'd6108;
        10'h2b2: pwm_thresh = 14'd6117;
        10'h2b3: pwm_thresh = 14'd6126;
        10'h2b4: pwm_thresh = 14'd6135;
        10'h2b5: pwm_thresh = 14'd6144;
        10'h2b6: pwm_thresh = 14'd6153;
        10'h2b7: pwm_thresh = 14'd6161;
        10'h2b8: pwm_thresh = 14'd6170;
        10'h2b9: pwm_thresh = 14'd6179;
        10'h2ba: pwm_thresh = 14'd6188;
        10'h2bb: pwm_thresh = 14'd6197;
        10'h2bc: pwm_thresh = 14'd6206;
        10'h2bd: pwm_thresh = 14'd6215;
        10'h2be: pwm_thresh = 14'd6223;
        10'h2bf: pwm_thresh = 14'd6232;
        10'h2c0: pwm_thresh = 14'd6241;
        10'h2c1: pwm_thresh = 14'd6250;
        10'h2c2: pwm_thresh = 14'd6259;
        10'h2c3: pwm_thresh = 14'd6268;
        10'h2c4: pwm_thresh = 14'd6277;
        10'h2c5: pwm_thresh = 14'd6286;
        10'h2c6: pwm_thresh = 14'd6294;
        10'h2c7: pwm_thresh = 14'd6303;
        10'h2c8: pwm_thresh = 14'd6312;
        10'h2c9: pwm_thresh = 14'd6321;
        10'h2ca: pwm_thresh = 14'd6330;
        10'h2cb: pwm_thresh = 14'd6339;
        10'h2cc: pwm_thresh = 14'd6348;
        10'h2cd: pwm_thresh = 14'd6356;
        10'h2ce: pwm_thresh = 14'd6365;
        10'h2cf: pwm_thresh = 14'd6374;
        10'h2d0: pwm_thresh = 14'd6383;
        10'h2d1: pwm_thresh = 14'd6392;
        10'h2d2: pwm_thresh = 14'd6401;
        10'h2d3: pwm_thresh = 14'd6410;
        10'h2d4: pwm_thresh = 14'd6419;
        10'h2d5: pwm_thresh = 14'd6427;
        10'h2d6: pwm_thresh = 14'd6436;
        10'h2d7: pwm_thresh = 14'd6445;
        10'h2d8: pwm_thresh = 14'd6454;
        10'h2d9: pwm_thresh = 14'd6463;
        10'h2da: pwm_thresh = 14'd6472;
        10'h2db: pwm_thresh = 14'd6481;
        10'h2dc: pwm_thresh = 14'd6489;
        10'h2dd: pwm_thresh = 14'd6498;
        10'h2de: pwm_thresh = 14'd6507;
        10'h2df: pwm_thresh = 14'd6516;
        10'h2e0: pwm_thresh = 14'd6525;
        10'h2e1: pwm_thresh = 14'd6534;
        10'h2e2: pwm_thresh = 14'd6543;
        10'h2e3: pwm_thresh = 14'd6552;
        10'h2e4: pwm_thresh = 14'd6560;
        10'h2e5: pwm_thresh = 14'd6569;
        10'h2e6: pwm_thresh = 14'd6578;
        10'h2e7: pwm_thresh = 14'd6587;
        10'h2e8: pwm_thresh = 14'd6596;
        10'h2e9: pwm_thresh = 14'd6605;
        10'h2ea: pwm_thresh = 14'd6614;
        10'h2eb: pwm_thresh = 14'd6622;
        10'h2ec: pwm_thresh = 14'd6631;
        10'h2ed: pwm_thresh = 14'd6640;
        10'h2ee: pwm_thresh = 14'd6649;
        10'h2ef: pwm_thresh = 14'd6658;
        10'h2f0: pwm_thresh = 14'd6667;
        10'h2f1: pwm_thresh = 14'd6676;
        10'h2f2: pwm_thresh = 14'd6685;
        10'h2f3: pwm_thresh = 14'd6693;
        10'h2f4: pwm_thresh = 14'd6702;
        10'h2f5: pwm_thresh = 14'd6711;
        10'h2f6: pwm_thresh = 14'd6720;
        10'h2f7: pwm_thresh = 14'd6729;
        10'h2f8: pwm_thresh = 14'd6738;
        10'h2f9: pwm_thresh = 14'd6747;
        10'h2fa: pwm_thresh = 14'd6755;
        10'h2fb: pwm_thresh = 14'd6764;
        10'h2fc: pwm_thresh = 14'd6773;
        10'h2fd: pwm_thresh = 14'd6782;
        10'h2fe: pwm_thresh = 14'd6791;
        10'h2ff: pwm_thresh = 14'd6800;
        10'h300: pwm_thresh = 14'd6809;
        10'h301: pwm_thresh = 14'd6818;
        10'h302: pwm_thresh = 14'd6826;
        10'h303: pwm_thresh = 14'd6835;
        10'h304: pwm_thresh = 14'd6844;
        10'h305: pwm_thresh = 14'd6853;
        10'h306: pwm_thresh = 14'd6862;
        10'h307: pwm_thresh = 14'd6871;
        10'h308: pwm_thresh = 14'd6880;
        10'h309: pwm_thresh = 14'd6888;
        10'h30a: pwm_thresh = 14'd6897;
        10'h30b: pwm_thresh = 14'd6906;
        10'h30c: pwm_thresh = 14'd6915;
        10'h30d: pwm_thresh = 14'd6924;
        10'h30e: pwm_thresh = 14'd6933;
        10'h30f: pwm_thresh = 14'd6942;
        10'h310: pwm_thresh = 14'd6951;
        10'h311: pwm_thresh = 14'd6959;
        10'h312: pwm_thresh = 14'd6968;
        10'h313: pwm_thresh = 14'd6977;
        10'h314: pwm_thresh = 14'd6986;
        10'h315: pwm_thresh = 14'd6995;
        10'h316: pwm_thresh = 14'd7004;
        10'h317: pwm_thresh = 14'd7013;
        10'h318: pwm_thresh = 14'd7021;
        10'h319: pwm_thresh = 14'd7030;
        10'h31a: pwm_thresh = 14'd7039;
        10'h31b: pwm_thresh = 14'd7048;
        10'h31c: pwm_thresh = 14'd7057;
        10'h31d: pwm_thresh = 14'd7066;
        10'h31e: pwm_thresh = 14'd7075;
        10'h31f: pwm_thresh = 14'd7083;
        10'h320: pwm_thresh = 14'd7092;
        10'h321: pwm_thresh = 14'd7101;
        10'h322: pwm_thresh = 14'd7110;
        10'h323: pwm_thresh = 14'd7119;
        10'h324: pwm_thresh = 14'd7128;
        10'h325: pwm_thresh = 14'd7137;
        10'h326: pwm_thresh = 14'd7146;
        10'h327: pwm_thresh = 14'd7154;
        10'h328: pwm_thresh = 14'd7163;
        10'h329: pwm_thresh = 14'd7172;
        10'h32a: pwm_thresh = 14'd7181;
        10'h32b: pwm_thresh = 14'd7190;
        10'h32c: pwm_thresh = 14'd7199;
        10'h32d: pwm_thresh = 14'd7208;
        10'h32e: pwm_thresh = 14'd7216;
        10'h32f: pwm_thresh = 14'd7225;
        10'h330: pwm_thresh = 14'd7234;
        10'h331: pwm_thresh = 14'd7243;
        10'h332: pwm_thresh = 14'd7252;
        10'h333: pwm_thresh = 14'd7261;
        10'h334: pwm_thresh = 14'd7270;
        10'h335: pwm_thresh = 14'd7279;
        10'h336: pwm_thresh = 14'd7287;
        10'h337: pwm_thresh = 14'd7296;
        10'h338: pwm_thresh = 14'd7305;
        10'h339: pwm_thresh = 14'd7314;
        10'h33a: pwm_thresh = 14'd7323;
        10'h33b: pwm_thresh = 14'd7332;
        10'h33c: pwm_thresh = 14'd7341;
        10'h33d: pwm_thresh = 14'd7349;
        10'h33e: pwm_thresh = 14'd7358;
        10'h33f: pwm_thresh = 14'd7367;
        10'h340: pwm_thresh = 14'd7376;
        10'h341: pwm_thresh = 14'd7385;
        10'h342: pwm_thresh = 14'd7394;
        10'h343: pwm_thresh = 14'd7403;
        10'h344: pwm_thresh = 14'd7412;
        10'h345: pwm_thresh = 14'd7420;
        10'h346: pwm_thresh = 14'd7429;
        10'h347: pwm_thresh = 14'd7438;
        10'h348: pwm_thresh = 14'd7447;
        10'h349: pwm_thresh = 14'd7456;
        10'h34a: pwm_thresh = 14'd7465;
        10'h34b: pwm_thresh = 14'd7474;
        10'h34c: pwm_thresh = 14'd7482;
        10'h34d: pwm_thresh = 14'd7491;
        10'h34e: pwm_thresh = 14'd7500;
        10'h34f: pwm_thresh = 14'd7509;
        10'h350: pwm_thresh = 14'd7518;
        10'h351: pwm_thresh = 14'd7527;
        10'h352: pwm_thresh = 14'd7536;
        10'h353: pwm_thresh = 14'd7545;
        10'h354: pwm_thresh = 14'd7553;
        10'h355: pwm_thresh = 14'd7562;
        10'h356: pwm_thresh = 14'd7571;
        10'h357: pwm_thresh = 14'd7580;
        10'h358: pwm_thresh = 14'd7589;
        10'h359: pwm_thresh = 14'd7598;
        10'h35a: pwm_thresh = 14'd7607;
        10'h35b: pwm_thresh = 14'd7615;
        10'h35c: pwm_thresh = 14'd7624;
        10'h35d: pwm_thresh = 14'd7633;
        10'h35e: pwm_thresh = 14'd7642;
        10'h35f: pwm_thresh = 14'd7651;
        10'h360: pwm_thresh = 14'd7660;
        10'h361: pwm_thresh = 14'd7669;
        10'h362: pwm_thresh = 14'd7678;
        10'h363: pwm_thresh = 14'd7686;
        10'h364: pwm_thresh = 14'd7695;
        10'h365: pwm_thresh = 14'd7704;
        10'h366: pwm_thresh = 14'd7713;
        10'h367: pwm_thresh = 14'd7722;
        10'h368: pwm_thresh = 14'd7731;
        10'h369: pwm_thresh = 14'd7740;
        10'h36a: pwm_thresh = 14'd7748;
        10'h36b: pwm_thresh = 14'd7757;
        10'h36c: pwm_thresh = 14'd7766;
        10'h36d: pwm_thresh = 14'd7775;
        10'h36e: pwm_thresh = 14'd7784;
        10'h36f: pwm_thresh = 14'd7793;
        10'h370: pwm_thresh = 14'd7802;
        10'h371: pwm_thresh = 14'd7811;
        10'h372: pwm_thresh = 14'd7819;
        10'h373: pwm_thresh = 14'd7828;
        10'h374: pwm_thresh = 14'd7837;
        10'h375: pwm_thresh = 14'd7846;
        10'h376: pwm_thresh = 14'd7855;
        10'h377: pwm_thresh = 14'd7864;
        10'h378: pwm_thresh = 14'd7873;
        10'h379: pwm_thresh = 14'd7881;
        10'h37a: pwm_thresh = 14'd7890;
        10'h37b: pwm_thresh = 14'd7899;
        10'h37c: pwm_thresh = 14'd7908;
        10'h37d: pwm_thresh = 14'd7917;
        10'h37e: pwm_thresh = 14'd7926;
        10'h37f: pwm_thresh = 14'd7935;
        10'h380: pwm_thresh = 14'd7944;
        10'h381: pwm_thresh = 14'd7952;
        10'h382: pwm_thresh = 14'd7961;
        10'h383: pwm_thresh = 14'd7970;
        10'h384: pwm_thresh = 14'd7979;
        10'h385: pwm_thresh = 14'd7988;
        10'h386: pwm_thresh = 14'd7997;
        10'h387: pwm_thresh = 14'd8006;
        10'h388: pwm_thresh = 14'd8014;
        10'h389: pwm_thresh = 14'd8023;
        10'h38a: pwm_thresh = 14'd8032;
        10'h38b: pwm_thresh = 14'd8041;
        10'h38c: pwm_thresh = 14'd8050;
        10'h38d: pwm_thresh = 14'd8059;
        10'h38e: pwm_thresh = 14'd8068;
        10'h38f: pwm_thresh = 14'd8076;
        10'h390: pwm_thresh = 14'd8085;
        10'h391: pwm_thresh = 14'd8094;
        10'h392: pwm_thresh = 14'd8103;
        10'h393: pwm_thresh = 14'd8112;
        10'h394: pwm_thresh = 14'd8121;
        10'h395: pwm_thresh = 14'd8130;
        10'h396: pwm_thresh = 14'd8139;
        10'h397: pwm_thresh = 14'd8147;
        10'h398: pwm_thresh = 14'd8156;
        10'h399: pwm_thresh = 14'd8165;
        10'h39a: pwm_thresh = 14'd8174;
        10'h39b: pwm_thresh = 14'd8183;
        10'h39c: pwm_thresh = 14'd8192;
        10'h39d: pwm_thresh = 14'd8201;
        10'h39e: pwm_thresh = 14'd8209;
        10'h39f: pwm_thresh = 14'd8218;
        10'h3a0: pwm_thresh = 14'd8227;
        10'h3a1: pwm_thresh = 14'd8236;
        10'h3a2: pwm_thresh = 14'd8245;
        10'h3a3: pwm_thresh = 14'd8254;
        10'h3a4: pwm_thresh = 14'd8263;
        10'h3a5: pwm_thresh = 14'd8272;
        10'h3a6: pwm_thresh = 14'd8280;
        10'h3a7: pwm_thresh = 14'd8289;
        10'h3a8: pwm_thresh = 14'd8298;
        10'h3a9: pwm_thresh = 14'd8307;
        10'h3aa: pwm_thresh = 14'd8316;
        10'h3ab: pwm_thresh = 14'd8325;
        10'h3ac: pwm_thresh = 14'd8334;
        10'h3ad: pwm_thresh = 14'd8342;
        10'h3ae: pwm_thresh = 14'd8351;
        10'h3af: pwm_thresh = 14'd8360;
        10'h3b0: pwm_thresh = 14'd8369;
        10'h3b1: pwm_thresh = 14'd8378;
        10'h3b2: pwm_thresh = 14'd8387;
        10'h3b3: pwm_thresh = 14'd8396;
        10'h3b4: pwm_thresh = 14'd8405;
        10'h3b5: pwm_thresh = 14'd8413;
        10'h3b6: pwm_thresh = 14'd8422;
        10'h3b7: pwm_thresh = 14'd8431;
        10'h3b8: pwm_thresh = 14'd8440;
        10'h3b9: pwm_thresh = 14'd8449;
        10'h3ba: pwm_thresh = 14'd8458;
        10'h3bb: pwm_thresh = 14'd8467;
        10'h3bc: pwm_thresh = 14'd8475;
        10'h3bd: pwm_thresh = 14'd8484;
        10'h3be: pwm_thresh = 14'd8493;
        10'h3bf: pwm_thresh = 14'd8502;
        10'h3c0: pwm_thresh = 14'd8511;
        10'h3c1: pwm_thresh = 14'd8520;
        10'h3c2: pwm_thresh = 14'd8529;
        10'h3c3: pwm_thresh = 14'd8538;
        10'h3c4: pwm_thresh = 14'd8546;
        10'h3c5: pwm_thresh = 14'd8555;
        10'h3c6: pwm_thresh = 14'd8564;
        10'h3c7: pwm_thresh = 14'd8573;
        10'h3c8: pwm_thresh = 14'd8582;
        10'h3c9: pwm_thresh = 14'd8591;
        10'h3ca: pwm_thresh = 14'd8600;
        10'h3cb: pwm_thresh = 14'd8608;
        10'h3cc: pwm_thresh = 14'd8617;
        10'h3cd: pwm_thresh = 14'd8626;
        10'h3ce: pwm_thresh = 14'd8635;
        10'h3cf: pwm_thresh = 14'd8644;
        10'h3d0: pwm_thresh = 14'd8653;
        10'h3d1: pwm_thresh = 14'd8662;
        10'h3d2: pwm_thresh = 14'd8671;
        10'h3d3: pwm_thresh = 14'd8679;
        10'h3d4: pwm_thresh = 14'd8688;
        10'h3d5: pwm_thresh = 14'd8697;
        10'h3d6: pwm_thresh = 14'd8706;
        10'h3d7: pwm_thresh = 14'd8715;
        10'h3d8: pwm_thresh = 14'd8724;
        10'h3d9: pwm_thresh = 14'd8733;
        10'h3da: pwm_thresh = 14'd8741;
        10'h3db: pwm_thresh = 14'd8750;
        10'h3dc: pwm_thresh = 14'd8759;
        10'h3dd: pwm_thresh = 14'd8768;
        10'h3de: pwm_thresh = 14'd8777;
        10'h3df: pwm_thresh = 14'd8786;
        10'h3e0: pwm_thresh = 14'd8795;
        10'h3e1: pwm_thresh = 14'd8804;
        10'h3e2: pwm_thresh = 14'd8812;
        10'h3e3: pwm_thresh = 14'd8821;
        10'h3e4: pwm_thresh = 14'd8830;
        10'h3e5: pwm_thresh = 14'd8839;
        10'h3e6: pwm_thresh = 14'd8848;
        10'h3e7: pwm_thresh = 14'd8857;
        10'h3e8: pwm_thresh = 14'd8866;
        10'h3e9: pwm_thresh = 14'd8874;
        10'h3ea: pwm_thresh = 14'd8883;
        10'h3eb: pwm_thresh = 14'd8892;
        10'h3ec: pwm_thresh = 14'd8901;
        10'h3ed: pwm_thresh = 14'd8910;
        10'h3ee: pwm_thresh = 14'd8919;
        10'h3ef: pwm_thresh = 14'd8928;
        10'h3f0: pwm_thresh = 14'd8937;
        10'h3f1: pwm_thresh = 14'd8945;
        10'h3f2: pwm_thresh = 14'd8954;
        10'h3f3: pwm_thresh = 14'd8963;
        10'h3f4: pwm_thresh = 14'd8972;
        10'h3f5: pwm_thresh = 14'd8981;
        10'h3f6: pwm_thresh = 14'd8990;
        10'h3f7: pwm_thresh = 14'd8999;
        10'h3f8: pwm_thresh = 14'd9007;
        10'h3f9: pwm_thresh = 14'd9016;
        10'h3fa: pwm_thresh = 14'd9025;
        10'h3fb: pwm_thresh = 14'd9034;
        10'h3fc: pwm_thresh = 14'd9043;
        10'h3fd: pwm_thresh = 14'd9052;
        10'h3fe: pwm_thresh = 14'd9061;
        10'h3ff: pwm_thresh = 14'd9070;
    endcase
  end

 
endmodule: pwm_thresh_father
