

module pwm_thresholder
  (input  logic [9:0] mult_val,
   output logic [26:0] pwm_thresh);

    always_comb begin
      case(mult_val)
      10'h0: pwm_thresh = 27'd0;
      10'h1: pwm_thresh = 27'd97751;
      10'h2: pwm_thresh = 27'd195503;
      10'h3: pwm_thresh = 27'd293255;
      10'h4: pwm_thresh = 27'd391006;
      10'h5: pwm_thresh = 27'd488758;
      10'h6: pwm_thresh = 27'd586510;
      10'h7: pwm_thresh = 27'd684261;
      10'h8: pwm_thresh = 27'd782013;
      10'h9: pwm_thresh = 27'd879765;
      10'ha: pwm_thresh = 27'd977517;
      10'hb: pwm_thresh = 27'd1075268;
      10'hc: pwm_thresh = 27'd1173020;
      10'hd: pwm_thresh = 27'd1270772;
      10'he: pwm_thresh = 27'd1368523;
      10'hf: pwm_thresh = 27'd1466275;
      10'h10: pwm_thresh = 27'd1564027;
      10'h11: pwm_thresh = 27'd1661779;
      10'h12: pwm_thresh = 27'd1759530;
      10'h13: pwm_thresh = 27'd1857282;
      10'h14: pwm_thresh = 27'd1955034;
      10'h15: pwm_thresh = 27'd2052785;
      10'h16: pwm_thresh = 27'd2150537;
      10'h17: pwm_thresh = 27'd2248289;
      10'h18: pwm_thresh = 27'd2346041;
      10'h19: pwm_thresh = 27'd2443792;
      10'h1a: pwm_thresh = 27'd2541544;
      10'h1b: pwm_thresh = 27'd2639296;
      10'h1c: pwm_thresh = 27'd2737047;
      10'h1d: pwm_thresh = 27'd2834799;
      10'h1e: pwm_thresh = 27'd2932551;
      10'h1f: pwm_thresh = 27'd3030303;
      10'h20: pwm_thresh = 27'd3128054;
      10'h21: pwm_thresh = 27'd3225806;
      10'h22: pwm_thresh = 27'd3323558;
      10'h23: pwm_thresh = 27'd3421309;
      10'h24: pwm_thresh = 27'd3519061;
      10'h25: pwm_thresh = 27'd3616813;
      10'h26: pwm_thresh = 27'd3714565;
      10'h27: pwm_thresh = 27'd3812316;
      10'h28: pwm_thresh = 27'd3910068;
      10'h29: pwm_thresh = 27'd4007820;
      10'h2a: pwm_thresh = 27'd4105571;
      10'h2b: pwm_thresh = 27'd4203323;
      10'h2c: pwm_thresh = 27'd4301075;
      10'h2d: pwm_thresh = 27'd4398826;
      10'h2e: pwm_thresh = 27'd4496578;
      10'h2f: pwm_thresh = 27'd4594330;
      10'h30: pwm_thresh = 27'd4692082;
      10'h31: pwm_thresh = 27'd4789833;
      10'h32: pwm_thresh = 27'd4887585;
      10'h33: pwm_thresh = 27'd4985337;
      10'h34: pwm_thresh = 27'd5083088;
      10'h35: pwm_thresh = 27'd5180840;
      10'h36: pwm_thresh = 27'd5278592;
      10'h37: pwm_thresh = 27'd5376344;
      10'h38: pwm_thresh = 27'd5474095;
      10'h39: pwm_thresh = 27'd5571847;
      10'h3a: pwm_thresh = 27'd5669599;
      10'h3b: pwm_thresh = 27'd5767350;
      10'h3c: pwm_thresh = 27'd5865102;
      10'h3d: pwm_thresh = 27'd5962854;
      10'h3e: pwm_thresh = 27'd6060606;
      10'h3f: pwm_thresh = 27'd6158357;
      10'h40: pwm_thresh = 27'd6256109;
      10'h41: pwm_thresh = 27'd6353861;
      10'h42: pwm_thresh = 27'd6451612;
      10'h43: pwm_thresh = 27'd6549364;
      10'h44: pwm_thresh = 27'd6647116;
      10'h45: pwm_thresh = 27'd6744868;
      10'h46: pwm_thresh = 27'd6842619;
      10'h47: pwm_thresh = 27'd6940371;
      10'h48: pwm_thresh = 27'd7038123;
      10'h49: pwm_thresh = 27'd7135874;
      10'h4a: pwm_thresh = 27'd7233626;
      10'h4b: pwm_thresh = 27'd7331378;
      10'h4c: pwm_thresh = 27'd7429130;
      10'h4d: pwm_thresh = 27'd7526881;
      10'h4e: pwm_thresh = 27'd7624633;
      10'h4f: pwm_thresh = 27'd7722385;
      10'h50: pwm_thresh = 27'd7820136;
      10'h51: pwm_thresh = 27'd7917888;
      10'h52: pwm_thresh = 27'd8015640;
      10'h53: pwm_thresh = 27'd8113391;
      10'h54: pwm_thresh = 27'd8211143;
      10'h55: pwm_thresh = 27'd8308895;
      10'h56: pwm_thresh = 27'd8406647;
      10'h57: pwm_thresh = 27'd8504398;
      10'h58: pwm_thresh = 27'd8602150;
      10'h59: pwm_thresh = 27'd8699902;
      10'h5a: pwm_thresh = 27'd8797653;
      10'h5b: pwm_thresh = 27'd8895405;
      10'h5c: pwm_thresh = 27'd8993157;
      10'h5d: pwm_thresh = 27'd9090909;
      10'h5e: pwm_thresh = 27'd9188660;
      10'h5f: pwm_thresh = 27'd9286412;
      10'h60: pwm_thresh = 27'd9384164;
      10'h61: pwm_thresh = 27'd9481915;
      10'h62: pwm_thresh = 27'd9579667;
      10'h63: pwm_thresh = 27'd9677419;
      10'h64: pwm_thresh = 27'd9775171;
      10'h65: pwm_thresh = 27'd9872922;
      10'h66: pwm_thresh = 27'd9970674;
      10'h67: pwm_thresh = 27'd10068426;
      10'h68: pwm_thresh = 27'd10166177;
      10'h69: pwm_thresh = 27'd10263929;
      10'h6a: pwm_thresh = 27'd10361681;
      10'h6b: pwm_thresh = 27'd10459433;
      10'h6c: pwm_thresh = 27'd10557184;
      10'h6d: pwm_thresh = 27'd10654936;
      10'h6e: pwm_thresh = 27'd10752688;
      10'h6f: pwm_thresh = 27'd10850439;
      10'h70: pwm_thresh = 27'd10948191;
      10'h71: pwm_thresh = 27'd11045943;
      10'h72: pwm_thresh = 27'd11143695;
      10'h73: pwm_thresh = 27'd11241446;
      10'h74: pwm_thresh = 27'd11339198;
      10'h75: pwm_thresh = 27'd11436950;
      10'h76: pwm_thresh = 27'd11534701;
      10'h77: pwm_thresh = 27'd11632453;
      10'h78: pwm_thresh = 27'd11730205;
      10'h79: pwm_thresh = 27'd11827956;
      10'h7a: pwm_thresh = 27'd11925708;
      10'h7b: pwm_thresh = 27'd12023460;
      10'h7c: pwm_thresh = 27'd12121212;
      10'h7d: pwm_thresh = 27'd12218963;
      10'h7e: pwm_thresh = 27'd12316715;
      10'h7f: pwm_thresh = 27'd12414467;
      10'h80: pwm_thresh = 27'd12512218;
      10'h81: pwm_thresh = 27'd12609970;
      10'h82: pwm_thresh = 27'd12707722;
      10'h83: pwm_thresh = 27'd12805474;
      10'h84: pwm_thresh = 27'd12903225;
      10'h85: pwm_thresh = 27'd13000977;
      10'h86: pwm_thresh = 27'd13098729;
      10'h87: pwm_thresh = 27'd13196480;
      10'h88: pwm_thresh = 27'd13294232;
      10'h89: pwm_thresh = 27'd13391984;
      10'h8a: pwm_thresh = 27'd13489736;
      10'h8b: pwm_thresh = 27'd13587487;
      10'h8c: pwm_thresh = 27'd13685239;
      10'h8d: pwm_thresh = 27'd13782991;
      10'h8e: pwm_thresh = 27'd13880742;
      10'h8f: pwm_thresh = 27'd13978494;
      10'h90: pwm_thresh = 27'd14076246;
      10'h91: pwm_thresh = 27'd14173998;
      10'h92: pwm_thresh = 27'd14271749;
      10'h93: pwm_thresh = 27'd14369501;
      10'h94: pwm_thresh = 27'd14467253;
      10'h95: pwm_thresh = 27'd14565004;
      10'h96: pwm_thresh = 27'd14662756;
      10'h97: pwm_thresh = 27'd14760508;
      10'h98: pwm_thresh = 27'd14858260;
      10'h99: pwm_thresh = 27'd14956011;
      10'h9a: pwm_thresh = 27'd15053763;
      10'h9b: pwm_thresh = 27'd15151515;
      10'h9c: pwm_thresh = 27'd15249266;
      10'h9d: pwm_thresh = 27'd15347018;
      10'h9e: pwm_thresh = 27'd15444770;
      10'h9f: pwm_thresh = 27'd15542521;
      10'ha0: pwm_thresh = 27'd15640273;
      10'ha1: pwm_thresh = 27'd15738025;
      10'ha2: pwm_thresh = 27'd15835777;
      10'ha3: pwm_thresh = 27'd15933528;
      10'ha4: pwm_thresh = 27'd16031280;
      10'ha5: pwm_thresh = 27'd16129032;
      10'ha6: pwm_thresh = 27'd16226783;
      10'ha7: pwm_thresh = 27'd16324535;
      10'ha8: pwm_thresh = 27'd16422287;
      10'ha9: pwm_thresh = 27'd16520039;
      10'haa: pwm_thresh = 27'd16617790;
      10'hab: pwm_thresh = 27'd16715542;
      10'hac: pwm_thresh = 27'd16813294;
      10'had: pwm_thresh = 27'd16911045;
      10'hae: pwm_thresh = 27'd17008797;
      10'haf: pwm_thresh = 27'd17106549;
      10'hb0: pwm_thresh = 27'd17204301;
      10'hb1: pwm_thresh = 27'd17302052;
      10'hb2: pwm_thresh = 27'd17399804;
      10'hb3: pwm_thresh = 27'd17497556;
      10'hb4: pwm_thresh = 27'd17595307;
      10'hb5: pwm_thresh = 27'd17693059;
      10'hb6: pwm_thresh = 27'd17790811;
      10'hb7: pwm_thresh = 27'd17888563;
      10'hb8: pwm_thresh = 27'd17986314;
      10'hb9: pwm_thresh = 27'd18084066;
      10'hba: pwm_thresh = 27'd18181818;
      10'hbb: pwm_thresh = 27'd18279569;
      10'hbc: pwm_thresh = 27'd18377321;
      10'hbd: pwm_thresh = 27'd18475073;
      10'hbe: pwm_thresh = 27'd18572825;
      10'hbf: pwm_thresh = 27'd18670576;
      10'hc0: pwm_thresh = 27'd18768328;
      10'hc1: pwm_thresh = 27'd18866080;
      10'hc2: pwm_thresh = 27'd18963831;
      10'hc3: pwm_thresh = 27'd19061583;
      10'hc4: pwm_thresh = 27'd19159335;
      10'hc5: pwm_thresh = 27'd19257086;
      10'hc6: pwm_thresh = 27'd19354838;
      10'hc7: pwm_thresh = 27'd19452590;
      10'hc8: pwm_thresh = 27'd19550342;
      10'hc9: pwm_thresh = 27'd19648093;
      10'hca: pwm_thresh = 27'd19745845;
      10'hcb: pwm_thresh = 27'd19843597;
      10'hcc: pwm_thresh = 27'd19941348;
      10'hcd: pwm_thresh = 27'd20039100;
      10'hce: pwm_thresh = 27'd20136852;
      10'hcf: pwm_thresh = 27'd20234604;
      10'hd0: pwm_thresh = 27'd20332355;
      10'hd1: pwm_thresh = 27'd20430107;
      10'hd2: pwm_thresh = 27'd20527859;
      10'hd3: pwm_thresh = 27'd20625610;
      10'hd4: pwm_thresh = 27'd20723362;
      10'hd5: pwm_thresh = 27'd20821114;
      10'hd6: pwm_thresh = 27'd20918866;
      10'hd7: pwm_thresh = 27'd21016617;
      10'hd8: pwm_thresh = 27'd21114369;
      10'hd9: pwm_thresh = 27'd21212121;
      10'hda: pwm_thresh = 27'd21309872;
      10'hdb: pwm_thresh = 27'd21407624;
      10'hdc: pwm_thresh = 27'd21505376;
      10'hdd: pwm_thresh = 27'd21603128;
      10'hde: pwm_thresh = 27'd21700879;
      10'hdf: pwm_thresh = 27'd21798631;
      10'he0: pwm_thresh = 27'd21896383;
      10'he1: pwm_thresh = 27'd21994134;
      10'he2: pwm_thresh = 27'd22091886;
      10'he3: pwm_thresh = 27'd22189638;
      10'he4: pwm_thresh = 27'd22287390;
      10'he5: pwm_thresh = 27'd22385141;
      10'he6: pwm_thresh = 27'd22482893;
      10'he7: pwm_thresh = 27'd22580645;
      10'he8: pwm_thresh = 27'd22678396;
      10'he9: pwm_thresh = 27'd22776148;
      10'hea: pwm_thresh = 27'd22873900;
      10'heb: pwm_thresh = 27'd22971652;
      10'hec: pwm_thresh = 27'd23069403;
      10'hed: pwm_thresh = 27'd23167155;
      10'hee: pwm_thresh = 27'd23264907;
      10'hef: pwm_thresh = 27'd23362658;
      10'hf0: pwm_thresh = 27'd23460410;
      10'hf1: pwm_thresh = 27'd23558162;
      10'hf2: pwm_thresh = 27'd23655913;
      10'hf3: pwm_thresh = 27'd23753665;
      10'hf4: pwm_thresh = 27'd23851417;
      10'hf5: pwm_thresh = 27'd23949169;
      10'hf6: pwm_thresh = 27'd24046920;
      10'hf7: pwm_thresh = 27'd24144672;
      10'hf8: pwm_thresh = 27'd24242424;
      10'hf9: pwm_thresh = 27'd24340175;
      10'hfa: pwm_thresh = 27'd24437927;
      10'hfb: pwm_thresh = 27'd24535679;
      10'hfc: pwm_thresh = 27'd24633431;
      10'hfd: pwm_thresh = 27'd24731182;
      10'hfe: pwm_thresh = 27'd24828934;
      10'hff: pwm_thresh = 27'd24926686;
      10'h100: pwm_thresh = 27'd25024437;
      10'h101: pwm_thresh = 27'd25122189;
      10'h102: pwm_thresh = 27'd25219941;
      10'h103: pwm_thresh = 27'd25317693;
      10'h104: pwm_thresh = 27'd25415444;
      10'h105: pwm_thresh = 27'd25513196;
      10'h106: pwm_thresh = 27'd25610948;
      10'h107: pwm_thresh = 27'd25708699;
      10'h108: pwm_thresh = 27'd25806451;
      10'h109: pwm_thresh = 27'd25904203;
      10'h10a: pwm_thresh = 27'd26001955;
      10'h10b: pwm_thresh = 27'd26099706;
      10'h10c: pwm_thresh = 27'd26197458;
      10'h10d: pwm_thresh = 27'd26295210;
      10'h10e: pwm_thresh = 27'd26392961;
      10'h10f: pwm_thresh = 27'd26490713;
      10'h110: pwm_thresh = 27'd26588465;
      10'h111: pwm_thresh = 27'd26686217;
      10'h112: pwm_thresh = 27'd26783968;
      10'h113: pwm_thresh = 27'd26881720;
      10'h114: pwm_thresh = 27'd26979472;
      10'h115: pwm_thresh = 27'd27077223;
      10'h116: pwm_thresh = 27'd27174975;
      10'h117: pwm_thresh = 27'd27272727;
      10'h118: pwm_thresh = 27'd27370478;
      10'h119: pwm_thresh = 27'd27468230;
      10'h11a: pwm_thresh = 27'd27565982;
      10'h11b: pwm_thresh = 27'd27663734;
      10'h11c: pwm_thresh = 27'd27761485;
      10'h11d: pwm_thresh = 27'd27859237;
      10'h11e: pwm_thresh = 27'd27956989;
      10'h11f: pwm_thresh = 27'd28054740;
      10'h120: pwm_thresh = 27'd28152492;
      10'h121: pwm_thresh = 27'd28250244;
      10'h122: pwm_thresh = 27'd28347996;
      10'h123: pwm_thresh = 27'd28445747;
      10'h124: pwm_thresh = 27'd28543499;
      10'h125: pwm_thresh = 27'd28641251;
      10'h126: pwm_thresh = 27'd28739002;
      10'h127: pwm_thresh = 27'd28836754;
      10'h128: pwm_thresh = 27'd28934506;
      10'h129: pwm_thresh = 27'd29032258;
      10'h12a: pwm_thresh = 27'd29130009;
      10'h12b: pwm_thresh = 27'd29227761;
      10'h12c: pwm_thresh = 27'd29325513;
      10'h12d: pwm_thresh = 27'd29423264;
      10'h12e: pwm_thresh = 27'd29521016;
      10'h12f: pwm_thresh = 27'd29618768;
      10'h130: pwm_thresh = 27'd29716520;
      10'h131: pwm_thresh = 27'd29814271;
      10'h132: pwm_thresh = 27'd29912023;
      10'h133: pwm_thresh = 27'd30009775;
      10'h134: pwm_thresh = 27'd30107526;
      10'h135: pwm_thresh = 27'd30205278;
      10'h136: pwm_thresh = 27'd30303030;
      10'h137: pwm_thresh = 27'd30400782;
      10'h138: pwm_thresh = 27'd30498533;
      10'h139: pwm_thresh = 27'd30596285;
      10'h13a: pwm_thresh = 27'd30694037;
      10'h13b: pwm_thresh = 27'd30791788;
      10'h13c: pwm_thresh = 27'd30889540;
      10'h13d: pwm_thresh = 27'd30987292;
      10'h13e: pwm_thresh = 27'd31085043;
      10'h13f: pwm_thresh = 27'd31182795;
      10'h140: pwm_thresh = 27'd31280547;
      10'h141: pwm_thresh = 27'd31378299;
      10'h142: pwm_thresh = 27'd31476050;
      10'h143: pwm_thresh = 27'd31573802;
      10'h144: pwm_thresh = 27'd31671554;
      10'h145: pwm_thresh = 27'd31769305;
      10'h146: pwm_thresh = 27'd31867057;
      10'h147: pwm_thresh = 27'd31964809;
      10'h148: pwm_thresh = 27'd32062561;
      10'h149: pwm_thresh = 27'd32160312;
      10'h14a: pwm_thresh = 27'd32258064;
      10'h14b: pwm_thresh = 27'd32355816;
      10'h14c: pwm_thresh = 27'd32453567;
      10'h14d: pwm_thresh = 27'd32551319;
      10'h14e: pwm_thresh = 27'd32649071;
      10'h14f: pwm_thresh = 27'd32746823;
      10'h150: pwm_thresh = 27'd32844574;
      10'h151: pwm_thresh = 27'd32942326;
      10'h152: pwm_thresh = 27'd33040078;
      10'h153: pwm_thresh = 27'd33137829;
      10'h154: pwm_thresh = 27'd33235581;
      10'h155: pwm_thresh = 27'd33333333;
      10'h156: pwm_thresh = 27'd33431085;
      10'h157: pwm_thresh = 27'd33528836;
      10'h158: pwm_thresh = 27'd33626588;
      10'h159: pwm_thresh = 27'd33724340;
      10'h15a: pwm_thresh = 27'd33822091;
      10'h15b: pwm_thresh = 27'd33919843;
      10'h15c: pwm_thresh = 27'd34017595;
      10'h15d: pwm_thresh = 27'd34115347;
      10'h15e: pwm_thresh = 27'd34213098;
      10'h15f: pwm_thresh = 27'd34310850;
      10'h160: pwm_thresh = 27'd34408602;
      10'h161: pwm_thresh = 27'd34506353;
      10'h162: pwm_thresh = 27'd34604105;
      10'h163: pwm_thresh = 27'd34701857;
      10'h164: pwm_thresh = 27'd34799608;
      10'h165: pwm_thresh = 27'd34897360;
      10'h166: pwm_thresh = 27'd34995112;
      10'h167: pwm_thresh = 27'd35092864;
      10'h168: pwm_thresh = 27'd35190615;
      10'h169: pwm_thresh = 27'd35288367;
      10'h16a: pwm_thresh = 27'd35386119;
      10'h16b: pwm_thresh = 27'd35483870;
      10'h16c: pwm_thresh = 27'd35581622;
      10'h16d: pwm_thresh = 27'd35679374;
      10'h16e: pwm_thresh = 27'd35777126;
      10'h16f: pwm_thresh = 27'd35874877;
      10'h170: pwm_thresh = 27'd35972629;
      10'h171: pwm_thresh = 27'd36070381;
      10'h172: pwm_thresh = 27'd36168132;
      10'h173: pwm_thresh = 27'd36265884;
      10'h174: pwm_thresh = 27'd36363636;
      10'h175: pwm_thresh = 27'd36461388;
      10'h176: pwm_thresh = 27'd36559139;
      10'h177: pwm_thresh = 27'd36656891;
      10'h178: pwm_thresh = 27'd36754643;
      10'h179: pwm_thresh = 27'd36852394;
      10'h17a: pwm_thresh = 27'd36950146;
      10'h17b: pwm_thresh = 27'd37047898;
      10'h17c: pwm_thresh = 27'd37145650;
      10'h17d: pwm_thresh = 27'd37243401;
      10'h17e: pwm_thresh = 27'd37341153;
      10'h17f: pwm_thresh = 27'd37438905;
      10'h180: pwm_thresh = 27'd37536656;
      10'h181: pwm_thresh = 27'd37634408;
      10'h182: pwm_thresh = 27'd37732160;
      10'h183: pwm_thresh = 27'd37829912;
      10'h184: pwm_thresh = 27'd37927663;
      10'h185: pwm_thresh = 27'd38025415;
      10'h186: pwm_thresh = 27'd38123167;
      10'h187: pwm_thresh = 27'd38220918;
      10'h188: pwm_thresh = 27'd38318670;
      10'h189: pwm_thresh = 27'd38416422;
      10'h18a: pwm_thresh = 27'd38514173;
      10'h18b: pwm_thresh = 27'd38611925;
      10'h18c: pwm_thresh = 27'd38709677;
      10'h18d: pwm_thresh = 27'd38807429;
      10'h18e: pwm_thresh = 27'd38905180;
      10'h18f: pwm_thresh = 27'd39002932;
      10'h190: pwm_thresh = 27'd39100684;
      10'h191: pwm_thresh = 27'd39198435;
      10'h192: pwm_thresh = 27'd39296187;
      10'h193: pwm_thresh = 27'd39393939;
      10'h194: pwm_thresh = 27'd39491691;
      10'h195: pwm_thresh = 27'd39589442;
      10'h196: pwm_thresh = 27'd39687194;
      10'h197: pwm_thresh = 27'd39784946;
      10'h198: pwm_thresh = 27'd39882697;
      10'h199: pwm_thresh = 27'd39980449;
      10'h19a: pwm_thresh = 27'd40078201;
      10'h19b: pwm_thresh = 27'd40175953;
      10'h19c: pwm_thresh = 27'd40273704;
      10'h19d: pwm_thresh = 27'd40371456;
      10'h19e: pwm_thresh = 27'd40469208;
      10'h19f: pwm_thresh = 27'd40566959;
      10'h1a0: pwm_thresh = 27'd40664711;
      10'h1a1: pwm_thresh = 27'd40762463;
      10'h1a2: pwm_thresh = 27'd40860215;
      10'h1a3: pwm_thresh = 27'd40957966;
      10'h1a4: pwm_thresh = 27'd41055718;
      10'h1a5: pwm_thresh = 27'd41153470;
      10'h1a6: pwm_thresh = 27'd41251221;
      10'h1a7: pwm_thresh = 27'd41348973;
      10'h1a8: pwm_thresh = 27'd41446725;
      10'h1a9: pwm_thresh = 27'd41544477;
      10'h1aa: pwm_thresh = 27'd41642228;
      10'h1ab: pwm_thresh = 27'd41739980;
      10'h1ac: pwm_thresh = 27'd41837732;
      10'h1ad: pwm_thresh = 27'd41935483;
      10'h1ae: pwm_thresh = 27'd42033235;
      10'h1af: pwm_thresh = 27'd42130987;
      10'h1b0: pwm_thresh = 27'd42228739;
      10'h1b1: pwm_thresh = 27'd42326490;
      10'h1b2: pwm_thresh = 27'd42424242;
      10'h1b3: pwm_thresh = 27'd42521994;
      10'h1b4: pwm_thresh = 27'd42619745;
      10'h1b5: pwm_thresh = 27'd42717497;
      10'h1b6: pwm_thresh = 27'd42815249;
      10'h1b7: pwm_thresh = 27'd42913000;
      10'h1b8: pwm_thresh = 27'd43010752;
      10'h1b9: pwm_thresh = 27'd43108504;
      10'h1ba: pwm_thresh = 27'd43206256;
      10'h1bb: pwm_thresh = 27'd43304007;
      10'h1bc: pwm_thresh = 27'd43401759;
      10'h1bd: pwm_thresh = 27'd43499511;
      10'h1be: pwm_thresh = 27'd43597262;
      10'h1bf: pwm_thresh = 27'd43695014;
      10'h1c0: pwm_thresh = 27'd43792766;
      10'h1c1: pwm_thresh = 27'd43890518;
      10'h1c2: pwm_thresh = 27'd43988269;
      10'h1c3: pwm_thresh = 27'd44086021;
      10'h1c4: pwm_thresh = 27'd44183773;
      10'h1c5: pwm_thresh = 27'd44281524;
      10'h1c6: pwm_thresh = 27'd44379276;
      10'h1c7: pwm_thresh = 27'd44477028;
      10'h1c8: pwm_thresh = 27'd44574780;
      10'h1c9: pwm_thresh = 27'd44672531;
      10'h1ca: pwm_thresh = 27'd44770283;
      10'h1cb: pwm_thresh = 27'd44868035;
      10'h1cc: pwm_thresh = 27'd44965786;
      10'h1cd: pwm_thresh = 27'd45063538;
      10'h1ce: pwm_thresh = 27'd45161290;
      10'h1cf: pwm_thresh = 27'd45259042;
      10'h1d0: pwm_thresh = 27'd45356793;
      10'h1d1: pwm_thresh = 27'd45454545;
      10'h1d2: pwm_thresh = 27'd45552297;
      10'h1d3: pwm_thresh = 27'd45650048;
      10'h1d4: pwm_thresh = 27'd45747800;
      10'h1d5: pwm_thresh = 27'd45845552;
      10'h1d6: pwm_thresh = 27'd45943304;
      10'h1d7: pwm_thresh = 27'd46041055;
      10'h1d8: pwm_thresh = 27'd46138807;
      10'h1d9: pwm_thresh = 27'd46236559;
      10'h1da: pwm_thresh = 27'd46334310;
      10'h1db: pwm_thresh = 27'd46432062;
      10'h1dc: pwm_thresh = 27'd46529814;
      10'h1dd: pwm_thresh = 27'd46627565;
      10'h1de: pwm_thresh = 27'd46725317;
      10'h1df: pwm_thresh = 27'd46823069;
      10'h1e0: pwm_thresh = 27'd46920821;
      10'h1e1: pwm_thresh = 27'd47018572;
      10'h1e2: pwm_thresh = 27'd47116324;
      10'h1e3: pwm_thresh = 27'd47214076;
      10'h1e4: pwm_thresh = 27'd47311827;
      10'h1e5: pwm_thresh = 27'd47409579;
      10'h1e6: pwm_thresh = 27'd47507331;
      10'h1e7: pwm_thresh = 27'd47605083;
      10'h1e8: pwm_thresh = 27'd47702834;
      10'h1e9: pwm_thresh = 27'd47800586;
      10'h1ea: pwm_thresh = 27'd47898338;
      10'h1eb: pwm_thresh = 27'd47996089;
      10'h1ec: pwm_thresh = 27'd48093841;
      10'h1ed: pwm_thresh = 27'd48191593;
      10'h1ee: pwm_thresh = 27'd48289345;
      10'h1ef: pwm_thresh = 27'd48387096;
      10'h1f0: pwm_thresh = 27'd48484848;
      10'h1f1: pwm_thresh = 27'd48582600;
      10'h1f2: pwm_thresh = 27'd48680351;
      10'h1f3: pwm_thresh = 27'd48778103;
      10'h1f4: pwm_thresh = 27'd48875855;
      10'h1f5: pwm_thresh = 27'd48973607;
      10'h1f6: pwm_thresh = 27'd49071358;
      10'h1f7: pwm_thresh = 27'd49169110;
      10'h1f8: pwm_thresh = 27'd49266862;
      10'h1f9: pwm_thresh = 27'd49364613;
      10'h1fa: pwm_thresh = 27'd49462365;
      10'h1fb: pwm_thresh = 27'd49560117;
      10'h1fc: pwm_thresh = 27'd49657869;
      10'h1fd: pwm_thresh = 27'd49755620;
      10'h1fe: pwm_thresh = 27'd49853372;
      10'h1ff: pwm_thresh = 27'd49951124;
      10'h200: pwm_thresh = 27'd50048875;
      10'h201: pwm_thresh = 27'd50146627;
      10'h202: pwm_thresh = 27'd50244379;
      10'h203: pwm_thresh = 27'd50342130;
      10'h204: pwm_thresh = 27'd50439882;
      10'h205: pwm_thresh = 27'd50537634;
      10'h206: pwm_thresh = 27'd50635386;
      10'h207: pwm_thresh = 27'd50733137;
      10'h208: pwm_thresh = 27'd50830889;
      10'h209: pwm_thresh = 27'd50928641;
      10'h20a: pwm_thresh = 27'd51026392;
      10'h20b: pwm_thresh = 27'd51124144;
      10'h20c: pwm_thresh = 27'd51221896;
      10'h20d: pwm_thresh = 27'd51319648;
      10'h20e: pwm_thresh = 27'd51417399;
      10'h20f: pwm_thresh = 27'd51515151;
      10'h210: pwm_thresh = 27'd51612903;
      10'h211: pwm_thresh = 27'd51710654;
      10'h212: pwm_thresh = 27'd51808406;
      10'h213: pwm_thresh = 27'd51906158;
      10'h214: pwm_thresh = 27'd52003910;
      10'h215: pwm_thresh = 27'd52101661;
      10'h216: pwm_thresh = 27'd52199413;
      10'h217: pwm_thresh = 27'd52297165;
      10'h218: pwm_thresh = 27'd52394916;
      10'h219: pwm_thresh = 27'd52492668;
      10'h21a: pwm_thresh = 27'd52590420;
      10'h21b: pwm_thresh = 27'd52688172;
      10'h21c: pwm_thresh = 27'd52785923;
      10'h21d: pwm_thresh = 27'd52883675;
      10'h21e: pwm_thresh = 27'd52981427;
      10'h21f: pwm_thresh = 27'd53079178;
      10'h220: pwm_thresh = 27'd53176930;
      10'h221: pwm_thresh = 27'd53274682;
      10'h222: pwm_thresh = 27'd53372434;
      10'h223: pwm_thresh = 27'd53470185;
      10'h224: pwm_thresh = 27'd53567937;
      10'h225: pwm_thresh = 27'd53665689;
      10'h226: pwm_thresh = 27'd53763440;
      10'h227: pwm_thresh = 27'd53861192;
      10'h228: pwm_thresh = 27'd53958944;
      10'h229: pwm_thresh = 27'd54056695;
      10'h22a: pwm_thresh = 27'd54154447;
      10'h22b: pwm_thresh = 27'd54252199;
      10'h22c: pwm_thresh = 27'd54349951;
      10'h22d: pwm_thresh = 27'd54447702;
      10'h22e: pwm_thresh = 27'd54545454;
      10'h22f: pwm_thresh = 27'd54643206;
      10'h230: pwm_thresh = 27'd54740957;
      10'h231: pwm_thresh = 27'd54838709;
      10'h232: pwm_thresh = 27'd54936461;
      10'h233: pwm_thresh = 27'd55034213;
      10'h234: pwm_thresh = 27'd55131964;
      10'h235: pwm_thresh = 27'd55229716;
      10'h236: pwm_thresh = 27'd55327468;
      10'h237: pwm_thresh = 27'd55425219;
      10'h238: pwm_thresh = 27'd55522971;
      10'h239: pwm_thresh = 27'd55620723;
      10'h23a: pwm_thresh = 27'd55718475;
      10'h23b: pwm_thresh = 27'd55816226;
      10'h23c: pwm_thresh = 27'd55913978;
      10'h23d: pwm_thresh = 27'd56011730;
      10'h23e: pwm_thresh = 27'd56109481;
      10'h23f: pwm_thresh = 27'd56207233;
      10'h240: pwm_thresh = 27'd56304985;
      10'h241: pwm_thresh = 27'd56402737;
      10'h242: pwm_thresh = 27'd56500488;
      10'h243: pwm_thresh = 27'd56598240;
      10'h244: pwm_thresh = 27'd56695992;
      10'h245: pwm_thresh = 27'd56793743;
      10'h246: pwm_thresh = 27'd56891495;
      10'h247: pwm_thresh = 27'd56989247;
      10'h248: pwm_thresh = 27'd57086999;
      10'h249: pwm_thresh = 27'd57184750;
      10'h24a: pwm_thresh = 27'd57282502;
      10'h24b: pwm_thresh = 27'd57380254;
      10'h24c: pwm_thresh = 27'd57478005;
      10'h24d: pwm_thresh = 27'd57575757;
      10'h24e: pwm_thresh = 27'd57673509;
      10'h24f: pwm_thresh = 27'd57771260;
      10'h250: pwm_thresh = 27'd57869012;
      10'h251: pwm_thresh = 27'd57966764;
      10'h252: pwm_thresh = 27'd58064516;
      10'h253: pwm_thresh = 27'd58162267;
      10'h254: pwm_thresh = 27'd58260019;
      10'h255: pwm_thresh = 27'd58357771;
      10'h256: pwm_thresh = 27'd58455522;
      10'h257: pwm_thresh = 27'd58553274;
      10'h258: pwm_thresh = 27'd58651026;
      10'h259: pwm_thresh = 27'd58748778;
      10'h25a: pwm_thresh = 27'd58846529;
      10'h25b: pwm_thresh = 27'd58944281;
      10'h25c: pwm_thresh = 27'd59042033;
      10'h25d: pwm_thresh = 27'd59139784;
      10'h25e: pwm_thresh = 27'd59237536;
      10'h25f: pwm_thresh = 27'd59335288;
      10'h260: pwm_thresh = 27'd59433040;
      10'h261: pwm_thresh = 27'd59530791;
      10'h262: pwm_thresh = 27'd59628543;
      10'h263: pwm_thresh = 27'd59726295;
      10'h264: pwm_thresh = 27'd59824046;
      10'h265: pwm_thresh = 27'd59921798;
      10'h266: pwm_thresh = 27'd60019550;
      10'h267: pwm_thresh = 27'd60117302;
      10'h268: pwm_thresh = 27'd60215053;
      10'h269: pwm_thresh = 27'd60312805;
      10'h26a: pwm_thresh = 27'd60410557;
      10'h26b: pwm_thresh = 27'd60508308;
      10'h26c: pwm_thresh = 27'd60606060;
      10'h26d: pwm_thresh = 27'd60703812;
      10'h26e: pwm_thresh = 27'd60801564;
      10'h26f: pwm_thresh = 27'd60899315;
      10'h270: pwm_thresh = 27'd60997067;
      10'h271: pwm_thresh = 27'd61094819;
      10'h272: pwm_thresh = 27'd61192570;
      10'h273: pwm_thresh = 27'd61290322;
      10'h274: pwm_thresh = 27'd61388074;
      10'h275: pwm_thresh = 27'd61485826;
      10'h276: pwm_thresh = 27'd61583577;
      10'h277: pwm_thresh = 27'd61681329;
      10'h278: pwm_thresh = 27'd61779081;
      10'h279: pwm_thresh = 27'd61876832;
      10'h27a: pwm_thresh = 27'd61974584;
      10'h27b: pwm_thresh = 27'd62072336;
      10'h27c: pwm_thresh = 27'd62170087;
      10'h27d: pwm_thresh = 27'd62267839;
      10'h27e: pwm_thresh = 27'd62365591;
      10'h27f: pwm_thresh = 27'd62463343;
      10'h280: pwm_thresh = 27'd62561094;
      10'h281: pwm_thresh = 27'd62658846;
      10'h282: pwm_thresh = 27'd62756598;
      10'h283: pwm_thresh = 27'd62854349;
      10'h284: pwm_thresh = 27'd62952101;
      10'h285: pwm_thresh = 27'd63049853;
      10'h286: pwm_thresh = 27'd63147605;
      10'h287: pwm_thresh = 27'd63245356;
      10'h288: pwm_thresh = 27'd63343108;
      10'h289: pwm_thresh = 27'd63440860;
      10'h28a: pwm_thresh = 27'd63538611;
      10'h28b: pwm_thresh = 27'd63636363;
      10'h28c: pwm_thresh = 27'd63734115;
      10'h28d: pwm_thresh = 27'd63831867;
      10'h28e: pwm_thresh = 27'd63929618;
      10'h28f: pwm_thresh = 27'd64027370;
      10'h290: pwm_thresh = 27'd64125122;
      10'h291: pwm_thresh = 27'd64222873;
      10'h292: pwm_thresh = 27'd64320625;
      10'h293: pwm_thresh = 27'd64418377;
      10'h294: pwm_thresh = 27'd64516129;
      10'h295: pwm_thresh = 27'd64613880;
      10'h296: pwm_thresh = 27'd64711632;
      10'h297: pwm_thresh = 27'd64809384;
      10'h298: pwm_thresh = 27'd64907135;
      10'h299: pwm_thresh = 27'd65004887;
      10'h29a: pwm_thresh = 27'd65102639;
      10'h29b: pwm_thresh = 27'd65200391;
      10'h29c: pwm_thresh = 27'd65298142;
      10'h29d: pwm_thresh = 27'd65395894;
      10'h29e: pwm_thresh = 27'd65493646;
      10'h29f: pwm_thresh = 27'd65591397;
      10'h2a0: pwm_thresh = 27'd65689149;
      10'h2a1: pwm_thresh = 27'd65786901;
      10'h2a2: pwm_thresh = 27'd65884652;
      10'h2a3: pwm_thresh = 27'd65982404;
      10'h2a4: pwm_thresh = 27'd66080156;
      10'h2a5: pwm_thresh = 27'd66177908;
      10'h2a6: pwm_thresh = 27'd66275659;
      10'h2a7: pwm_thresh = 27'd66373411;
      10'h2a8: pwm_thresh = 27'd66471163;
      10'h2a9: pwm_thresh = 27'd66568914;
      10'h2aa: pwm_thresh = 27'd66666666;
      10'h2ab: pwm_thresh = 27'd66764418;
      10'h2ac: pwm_thresh = 27'd66862170;
      10'h2ad: pwm_thresh = 27'd66959921;
      10'h2ae: pwm_thresh = 27'd67057673;
      10'h2af: pwm_thresh = 27'd67155425;
      10'h2b0: pwm_thresh = 27'd67253176;
      10'h2b1: pwm_thresh = 27'd67350928;
      10'h2b2: pwm_thresh = 27'd67448680;
      10'h2b3: pwm_thresh = 27'd67546432;
      10'h2b4: pwm_thresh = 27'd67644183;
      10'h2b5: pwm_thresh = 27'd67741935;
      10'h2b6: pwm_thresh = 27'd67839687;
      10'h2b7: pwm_thresh = 27'd67937438;
      10'h2b8: pwm_thresh = 27'd68035190;
      10'h2b9: pwm_thresh = 27'd68132942;
      10'h2ba: pwm_thresh = 27'd68230694;
      10'h2bb: pwm_thresh = 27'd68328445;
      10'h2bc: pwm_thresh = 27'd68426197;
      10'h2bd: pwm_thresh = 27'd68523949;
      10'h2be: pwm_thresh = 27'd68621700;
      10'h2bf: pwm_thresh = 27'd68719452;
      10'h2c0: pwm_thresh = 27'd68817204;
      10'h2c1: pwm_thresh = 27'd68914956;
      10'h2c2: pwm_thresh = 27'd69012707;
      10'h2c3: pwm_thresh = 27'd69110459;
      10'h2c4: pwm_thresh = 27'd69208211;
      10'h2c5: pwm_thresh = 27'd69305962;
      10'h2c6: pwm_thresh = 27'd69403714;
      10'h2c7: pwm_thresh = 27'd69501466;
      10'h2c8: pwm_thresh = 27'd69599217;
      10'h2c9: pwm_thresh = 27'd69696969;
      10'h2ca: pwm_thresh = 27'd69794721;
      10'h2cb: pwm_thresh = 27'd69892473;
      10'h2cc: pwm_thresh = 27'd69990224;
      10'h2cd: pwm_thresh = 27'd70087976;
      10'h2ce: pwm_thresh = 27'd70185728;
      10'h2cf: pwm_thresh = 27'd70283479;
      10'h2d0: pwm_thresh = 27'd70381231;
      10'h2d1: pwm_thresh = 27'd70478983;
      10'h2d2: pwm_thresh = 27'd70576735;
      10'h2d3: pwm_thresh = 27'd70674486;
      10'h2d4: pwm_thresh = 27'd70772238;
      10'h2d5: pwm_thresh = 27'd70869990;
      10'h2d6: pwm_thresh = 27'd70967741;
      10'h2d7: pwm_thresh = 27'd71065493;
      10'h2d8: pwm_thresh = 27'd71163245;
      10'h2d9: pwm_thresh = 27'd71260997;
      10'h2da: pwm_thresh = 27'd71358748;
      10'h2db: pwm_thresh = 27'd71456500;
      10'h2dc: pwm_thresh = 27'd71554252;
      10'h2dd: pwm_thresh = 27'd71652003;
      10'h2de: pwm_thresh = 27'd71749755;
      10'h2df: pwm_thresh = 27'd71847507;
      10'h2e0: pwm_thresh = 27'd71945259;
      10'h2e1: pwm_thresh = 27'd72043010;
      10'h2e2: pwm_thresh = 27'd72140762;
      10'h2e3: pwm_thresh = 27'd72238514;
      10'h2e4: pwm_thresh = 27'd72336265;
      10'h2e5: pwm_thresh = 27'd72434017;
      10'h2e6: pwm_thresh = 27'd72531769;
      10'h2e7: pwm_thresh = 27'd72629521;
      10'h2e8: pwm_thresh = 27'd72727272;
      10'h2e9: pwm_thresh = 27'd72825024;
      10'h2ea: pwm_thresh = 27'd72922776;
      10'h2eb: pwm_thresh = 27'd73020527;
      10'h2ec: pwm_thresh = 27'd73118279;
      10'h2ed: pwm_thresh = 27'd73216031;
      10'h2ee: pwm_thresh = 27'd73313782;
      10'h2ef: pwm_thresh = 27'd73411534;
      10'h2f0: pwm_thresh = 27'd73509286;
      10'h2f1: pwm_thresh = 27'd73607038;
      10'h2f2: pwm_thresh = 27'd73704789;
      10'h2f3: pwm_thresh = 27'd73802541;
      10'h2f4: pwm_thresh = 27'd73900293;
      10'h2f5: pwm_thresh = 27'd73998044;
      10'h2f6: pwm_thresh = 27'd74095796;
      10'h2f7: pwm_thresh = 27'd74193548;
      10'h2f8: pwm_thresh = 27'd74291300;
      10'h2f9: pwm_thresh = 27'd74389051;
      10'h2fa: pwm_thresh = 27'd74486803;
      10'h2fb: pwm_thresh = 27'd74584555;
      10'h2fc: pwm_thresh = 27'd74682306;
      10'h2fd: pwm_thresh = 27'd74780058;
      10'h2fe: pwm_thresh = 27'd74877810;
      10'h2ff: pwm_thresh = 27'd74975562;
      10'h300: pwm_thresh = 27'd75073313;
      10'h301: pwm_thresh = 27'd75171065;
      10'h302: pwm_thresh = 27'd75268817;
      10'h303: pwm_thresh = 27'd75366568;
      10'h304: pwm_thresh = 27'd75464320;
      10'h305: pwm_thresh = 27'd75562072;
      10'h306: pwm_thresh = 27'd75659824;
      10'h307: pwm_thresh = 27'd75757575;
      10'h308: pwm_thresh = 27'd75855327;
      10'h309: pwm_thresh = 27'd75953079;
      10'h30a: pwm_thresh = 27'd76050830;
      10'h30b: pwm_thresh = 27'd76148582;
      10'h30c: pwm_thresh = 27'd76246334;
      10'h30d: pwm_thresh = 27'd76344086;
      10'h30e: pwm_thresh = 27'd76441837;
      10'h30f: pwm_thresh = 27'd76539589;
      10'h310: pwm_thresh = 27'd76637341;
      10'h311: pwm_thresh = 27'd76735092;
      10'h312: pwm_thresh = 27'd76832844;
      10'h313: pwm_thresh = 27'd76930596;
      10'h314: pwm_thresh = 27'd77028347;
      10'h315: pwm_thresh = 27'd77126099;
      10'h316: pwm_thresh = 27'd77223851;
      10'h317: pwm_thresh = 27'd77321603;
      10'h318: pwm_thresh = 27'd77419354;
      10'h319: pwm_thresh = 27'd77517106;
      10'h31a: pwm_thresh = 27'd77614858;
      10'h31b: pwm_thresh = 27'd77712609;
      10'h31c: pwm_thresh = 27'd77810361;
      10'h31d: pwm_thresh = 27'd77908113;
      10'h31e: pwm_thresh = 27'd78005865;
      10'h31f: pwm_thresh = 27'd78103616;
      10'h320: pwm_thresh = 27'd78201368;
      10'h321: pwm_thresh = 27'd78299120;
      10'h322: pwm_thresh = 27'd78396871;
      10'h323: pwm_thresh = 27'd78494623;
      10'h324: pwm_thresh = 27'd78592375;
      10'h325: pwm_thresh = 27'd78690127;
      10'h326: pwm_thresh = 27'd78787878;
      10'h327: pwm_thresh = 27'd78885630;
      10'h328: pwm_thresh = 27'd78983382;
      10'h329: pwm_thresh = 27'd79081133;
      10'h32a: pwm_thresh = 27'd79178885;
      10'h32b: pwm_thresh = 27'd79276637;
      10'h32c: pwm_thresh = 27'd79374389;
      10'h32d: pwm_thresh = 27'd79472140;
      10'h32e: pwm_thresh = 27'd79569892;
      10'h32f: pwm_thresh = 27'd79667644;
      10'h330: pwm_thresh = 27'd79765395;
      10'h331: pwm_thresh = 27'd79863147;
      10'h332: pwm_thresh = 27'd79960899;
      10'h333: pwm_thresh = 27'd80058651;
      10'h334: pwm_thresh = 27'd80156402;
      10'h335: pwm_thresh = 27'd80254154;
      10'h336: pwm_thresh = 27'd80351906;
      10'h337: pwm_thresh = 27'd80449657;
      10'h338: pwm_thresh = 27'd80547409;
      10'h339: pwm_thresh = 27'd80645161;
      10'h33a: pwm_thresh = 27'd80742913;
      10'h33b: pwm_thresh = 27'd80840664;
      10'h33c: pwm_thresh = 27'd80938416;
      10'h33d: pwm_thresh = 27'd81036168;
      10'h33e: pwm_thresh = 27'd81133919;
      10'h33f: pwm_thresh = 27'd81231671;
      10'h340: pwm_thresh = 27'd81329423;
      10'h341: pwm_thresh = 27'd81427174;
      10'h342: pwm_thresh = 27'd81524926;
      10'h343: pwm_thresh = 27'd81622678;
      10'h344: pwm_thresh = 27'd81720430;
      10'h345: pwm_thresh = 27'd81818181;
      10'h346: pwm_thresh = 27'd81915933;
      10'h347: pwm_thresh = 27'd82013685;
      10'h348: pwm_thresh = 27'd82111436;
      10'h349: pwm_thresh = 27'd82209188;
      10'h34a: pwm_thresh = 27'd82306940;
      10'h34b: pwm_thresh = 27'd82404692;
      10'h34c: pwm_thresh = 27'd82502443;
      10'h34d: pwm_thresh = 27'd82600195;
      10'h34e: pwm_thresh = 27'd82697947;
      10'h34f: pwm_thresh = 27'd82795698;
      10'h350: pwm_thresh = 27'd82893450;
      10'h351: pwm_thresh = 27'd82991202;
      10'h352: pwm_thresh = 27'd83088954;
      10'h353: pwm_thresh = 27'd83186705;
      10'h354: pwm_thresh = 27'd83284457;
      10'h355: pwm_thresh = 27'd83382209;
      10'h356: pwm_thresh = 27'd83479960;
      10'h357: pwm_thresh = 27'd83577712;
      10'h358: pwm_thresh = 27'd83675464;
      10'h359: pwm_thresh = 27'd83773216;
      10'h35a: pwm_thresh = 27'd83870967;
      10'h35b: pwm_thresh = 27'd83968719;
      10'h35c: pwm_thresh = 27'd84066471;
      10'h35d: pwm_thresh = 27'd84164222;
      10'h35e: pwm_thresh = 27'd84261974;
      10'h35f: pwm_thresh = 27'd84359726;
      10'h360: pwm_thresh = 27'd84457478;
      10'h361: pwm_thresh = 27'd84555229;
      10'h362: pwm_thresh = 27'd84652981;
      10'h363: pwm_thresh = 27'd84750733;
      10'h364: pwm_thresh = 27'd84848484;
      10'h365: pwm_thresh = 27'd84946236;
      10'h366: pwm_thresh = 27'd85043988;
      10'h367: pwm_thresh = 27'd85141739;
      10'h368: pwm_thresh = 27'd85239491;
      10'h369: pwm_thresh = 27'd85337243;
      10'h36a: pwm_thresh = 27'd85434995;
      10'h36b: pwm_thresh = 27'd85532746;
      10'h36c: pwm_thresh = 27'd85630498;
      10'h36d: pwm_thresh = 27'd85728250;
      10'h36e: pwm_thresh = 27'd85826001;
      10'h36f: pwm_thresh = 27'd85923753;
      10'h370: pwm_thresh = 27'd86021505;
      10'h371: pwm_thresh = 27'd86119257;
      10'h372: pwm_thresh = 27'd86217008;
      10'h373: pwm_thresh = 27'd86314760;
      10'h374: pwm_thresh = 27'd86412512;
      10'h375: pwm_thresh = 27'd86510263;
      10'h376: pwm_thresh = 27'd86608015;
      10'h377: pwm_thresh = 27'd86705767;
      10'h378: pwm_thresh = 27'd86803519;
      10'h379: pwm_thresh = 27'd86901270;
      10'h37a: pwm_thresh = 27'd86999022;
      10'h37b: pwm_thresh = 27'd87096774;
      10'h37c: pwm_thresh = 27'd87194525;
      10'h37d: pwm_thresh = 27'd87292277;
      10'h37e: pwm_thresh = 27'd87390029;
      10'h37f: pwm_thresh = 27'd87487781;
      10'h380: pwm_thresh = 27'd87585532;
      10'h381: pwm_thresh = 27'd87683284;
      10'h382: pwm_thresh = 27'd87781036;
      10'h383: pwm_thresh = 27'd87878787;
      10'h384: pwm_thresh = 27'd87976539;
      10'h385: pwm_thresh = 27'd88074291;
      10'h386: pwm_thresh = 27'd88172043;
      10'h387: pwm_thresh = 27'd88269794;
      10'h388: pwm_thresh = 27'd88367546;
      10'h389: pwm_thresh = 27'd88465298;
      10'h38a: pwm_thresh = 27'd88563049;
      10'h38b: pwm_thresh = 27'd88660801;
      10'h38c: pwm_thresh = 27'd88758553;
      10'h38d: pwm_thresh = 27'd88856304;
      10'h38e: pwm_thresh = 27'd88954056;
      10'h38f: pwm_thresh = 27'd89051808;
      10'h390: pwm_thresh = 27'd89149560;
      10'h391: pwm_thresh = 27'd89247311;
      10'h392: pwm_thresh = 27'd89345063;
      10'h393: pwm_thresh = 27'd89442815;
      10'h394: pwm_thresh = 27'd89540566;
      10'h395: pwm_thresh = 27'd89638318;
      10'h396: pwm_thresh = 27'd89736070;
      10'h397: pwm_thresh = 27'd89833822;
      10'h398: pwm_thresh = 27'd89931573;
      10'h399: pwm_thresh = 27'd90029325;
      10'h39a: pwm_thresh = 27'd90127077;
      10'h39b: pwm_thresh = 27'd90224828;
      10'h39c: pwm_thresh = 27'd90322580;
      10'h39d: pwm_thresh = 27'd90420332;
      10'h39e: pwm_thresh = 27'd90518084;
      10'h39f: pwm_thresh = 27'd90615835;
      10'h3a0: pwm_thresh = 27'd90713587;
      10'h3a1: pwm_thresh = 27'd90811339;
      10'h3a2: pwm_thresh = 27'd90909090;
      10'h3a3: pwm_thresh = 27'd91006842;
      10'h3a4: pwm_thresh = 27'd91104594;
      10'h3a5: pwm_thresh = 27'd91202346;
      10'h3a6: pwm_thresh = 27'd91300097;
      10'h3a7: pwm_thresh = 27'd91397849;
      10'h3a8: pwm_thresh = 27'd91495601;
      10'h3a9: pwm_thresh = 27'd91593352;
      10'h3aa: pwm_thresh = 27'd91691104;
      10'h3ab: pwm_thresh = 27'd91788856;
      10'h3ac: pwm_thresh = 27'd91886608;
      10'h3ad: pwm_thresh = 27'd91984359;
      10'h3ae: pwm_thresh = 27'd92082111;
      10'h3af: pwm_thresh = 27'd92179863;
      10'h3b0: pwm_thresh = 27'd92277614;
      10'h3b1: pwm_thresh = 27'd92375366;
      10'h3b2: pwm_thresh = 27'd92473118;
      10'h3b3: pwm_thresh = 27'd92570869;
      10'h3b4: pwm_thresh = 27'd92668621;
      10'h3b5: pwm_thresh = 27'd92766373;
      10'h3b6: pwm_thresh = 27'd92864125;
      10'h3b7: pwm_thresh = 27'd92961876;
      10'h3b8: pwm_thresh = 27'd93059628;
      10'h3b9: pwm_thresh = 27'd93157380;
      10'h3ba: pwm_thresh = 27'd93255131;
      10'h3bb: pwm_thresh = 27'd93352883;
      10'h3bc: pwm_thresh = 27'd93450635;
      10'h3bd: pwm_thresh = 27'd93548387;
      10'h3be: pwm_thresh = 27'd93646138;
      10'h3bf: pwm_thresh = 27'd93743890;
      10'h3c0: pwm_thresh = 27'd93841642;
      10'h3c1: pwm_thresh = 27'd93939393;
      10'h3c2: pwm_thresh = 27'd94037145;
      10'h3c3: pwm_thresh = 27'd94134897;
      10'h3c4: pwm_thresh = 27'd94232649;
      10'h3c5: pwm_thresh = 27'd94330400;
      10'h3c6: pwm_thresh = 27'd94428152;
      10'h3c7: pwm_thresh = 27'd94525904;
      10'h3c8: pwm_thresh = 27'd94623655;
      10'h3c9: pwm_thresh = 27'd94721407;
      10'h3ca: pwm_thresh = 27'd94819159;
      10'h3cb: pwm_thresh = 27'd94916911;
      10'h3cc: pwm_thresh = 27'd95014662;
      10'h3cd: pwm_thresh = 27'd95112414;
      10'h3ce: pwm_thresh = 27'd95210166;
      10'h3cf: pwm_thresh = 27'd95307917;
      10'h3d0: pwm_thresh = 27'd95405669;
      10'h3d1: pwm_thresh = 27'd95503421;
      10'h3d2: pwm_thresh = 27'd95601173;
      10'h3d3: pwm_thresh = 27'd95698924;
      10'h3d4: pwm_thresh = 27'd95796676;
      10'h3d5: pwm_thresh = 27'd95894428;
      10'h3d6: pwm_thresh = 27'd95992179;
      10'h3d7: pwm_thresh = 27'd96089931;
      10'h3d8: pwm_thresh = 27'd96187683;
      10'h3d9: pwm_thresh = 27'd96285434;
      10'h3da: pwm_thresh = 27'd96383186;
      10'h3db: pwm_thresh = 27'd96480938;
      10'h3dc: pwm_thresh = 27'd96578690;
      10'h3dd: pwm_thresh = 27'd96676441;
      10'h3de: pwm_thresh = 27'd96774193;
      10'h3df: pwm_thresh = 27'd96871945;
      10'h3e0: pwm_thresh = 27'd96969696;
      10'h3e1: pwm_thresh = 27'd97067448;
      10'h3e2: pwm_thresh = 27'd97165200;
      10'h3e3: pwm_thresh = 27'd97262952;
      10'h3e4: pwm_thresh = 27'd97360703;
      10'h3e5: pwm_thresh = 27'd97458455;
      10'h3e6: pwm_thresh = 27'd97556207;
      10'h3e7: pwm_thresh = 27'd97653958;
      10'h3e8: pwm_thresh = 27'd97751710;
      10'h3e9: pwm_thresh = 27'd97849462;
      10'h3ea: pwm_thresh = 27'd97947214;
      10'h3eb: pwm_thresh = 27'd98044965;
      10'h3ec: pwm_thresh = 27'd98142717;
      10'h3ed: pwm_thresh = 27'd98240469;
      10'h3ee: pwm_thresh = 27'd98338220;
      10'h3ef: pwm_thresh = 27'd98435972;
      10'h3f0: pwm_thresh = 27'd98533724;
      10'h3f1: pwm_thresh = 27'd98631476;
      10'h3f2: pwm_thresh = 27'd98729227;
      10'h3f3: pwm_thresh = 27'd98826979;
      10'h3f4: pwm_thresh = 27'd98924731;
      10'h3f5: pwm_thresh = 27'd99022482;
      10'h3f6: pwm_thresh = 27'd99120234;
      10'h3f7: pwm_thresh = 27'd99217986;
      10'h3f8: pwm_thresh = 27'd99315738;
      10'h3f9: pwm_thresh = 27'd99413489;
      10'h3fa: pwm_thresh = 27'd99511241;
      10'h3fb: pwm_thresh = 27'd99608993;
      10'h3fc: pwm_thresh = 27'd99706744;
      10'h3fd: pwm_thresh = 27'd99804496;
      10'h3fe: pwm_thresh = 27'd99902248;
      10'h3ff: pwm_thresh = 27'd100000000;
      endcase
    end

endmodule: pwm_thresholder
